(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h46b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire0;
  input wire signed [(4'ha):(1'h0)] wire1;
  input wire signed [(5'h14):(1'h0)] wire2;
  input wire [(4'hf):(1'h0)] wire3;
  input wire signed [(5'h10):(1'h0)] wire4;
  wire [(5'h11):(1'h0)] wire970;
  wire [(4'hf):(1'h0)] wire470;
  wire signed [(3'h5):(1'h0)] wire468;
  wire [(5'h16):(1'h0)] wire310;
  wire signed [(5'h15):(1'h0)] wire5;
  wire signed [(3'h6):(1'h0)] wire33;
  wire [(5'h17):(1'h0)] wire34;
  wire signed [(5'h17):(1'h0)] wire35;
  wire signed [(4'ha):(1'h0)] wire308;
  reg [(5'h18):(1'h0)] reg351 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg350 = (1'h0);
  reg [(4'he):(1'h0)] reg348 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg347 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg346 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg345 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg343 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg342 = (1'h0);
  reg [(3'h5):(1'h0)] reg339 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg337 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg335 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg333 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg331 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg330 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg329 = (1'h0);
  reg [(4'ha):(1'h0)] reg328 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg319 = (1'h0);
  reg [(3'h5):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg316 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg315 = (1'h0);
  reg [(5'h10):(1'h0)] reg312 = (1'h0);
  reg [(5'h16):(1'h0)] reg311 = (1'h0);
  reg [(3'h4):(1'h0)] reg31 = (1'h0);
  reg [(5'h17):(1'h0)] reg30 = (1'h0);
  reg [(5'h14):(1'h0)] reg29 = (1'h0);
  reg [(2'h3):(1'h0)] reg27 = (1'h0);
  reg [(5'h15):(1'h0)] reg25 = (1'h0);
  reg [(5'h16):(1'h0)] reg24 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg18 = (1'h0);
  reg [(5'h18):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg14 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg13 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg10 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg9 = (1'h0);
  reg [(5'h12):(1'h0)] reg471 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg474 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg475 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg473 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg472 = (1'h0);
  reg [(3'h7):(1'h0)] reg352 = (1'h0);
  reg [(5'h14):(1'h0)] reg349 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg344 = (1'h0);
  reg [(4'hf):(1'h0)] reg341 = (1'h0);
  reg [(4'hb):(1'h0)] reg340 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg338 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg336 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg334 = (1'h0);
  reg [(4'ha):(1'h0)] forvar331 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg332 = (1'h0);
  reg [(5'h16):(1'h0)] reg327 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar326 = (1'h0);
  reg [(4'hf):(1'h0)] reg325 = (1'h0);
  reg [(2'h2):(1'h0)] reg324 = (1'h0);
  reg [(5'h11):(1'h0)] reg323 = (1'h0);
  reg [(5'h17):(1'h0)] forvar321 = (1'h0);
  reg [(5'h13):(1'h0)] forvar320 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg314 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg313 = (1'h0);
  reg [(5'h11):(1'h0)] forvar312 = (1'h0);
  reg signed [(4'he):(1'h0)] reg32 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg28 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar26 = (1'h0);
  reg [(2'h3):(1'h0)] reg23 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar22 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg21 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar12 = (1'h0);
  reg [(3'h4):(1'h0)] reg19 = (1'h0);
  reg [(4'hb):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg12 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg11 = (1'h0);
  reg [(4'h9):(1'h0)] reg8 = (1'h0);
  reg [(2'h2):(1'h0)] forvar7 = (1'h0);
  reg [(4'hd):(1'h0)] reg6 = (1'h0);
  assign y = {wire970,
                 wire470,
                 wire468,
                 wire310,
                 wire5,
                 wire33,
                 wire34,
                 wire35,
                 wire308,
                 reg351,
                 reg350,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg343,
                 reg342,
                 reg339,
                 reg337,
                 reg335,
                 reg333,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg322,
                 reg319,
                 reg318,
                 reg316,
                 reg315,
                 reg312,
                 reg311,
                 reg31,
                 reg30,
                 reg29,
                 reg27,
                 reg25,
                 reg24,
                 reg20,
                 reg18,
                 reg16,
                 reg14,
                 reg13,
                 reg10,
                 reg9,
                 reg471,
                 reg474,
                 reg475,
                 reg473,
                 reg472,
                 reg352,
                 reg349,
                 reg344,
                 reg341,
                 reg340,
                 reg338,
                 reg336,
                 reg334,
                 forvar331,
                 reg332,
                 reg327,
                 forvar326,
                 reg325,
                 reg324,
                 reg323,
                 forvar321,
                 forvar320,
                 reg317,
                 reg314,
                 reg313,
                 forvar312,
                 reg32,
                 reg28,
                 forvar26,
                 reg23,
                 forvar22,
                 reg21,
                 forvar12,
                 reg19,
                 reg17,
                 reg15,
                 reg12,
                 reg11,
                 reg8,
                 forvar7,
                 reg6,
                 (1'h0)};
  assign wire5 = (({(~|wire4[(4'h9):(2'h3)])} ?
                     (wire3 ?
                         ((wire0 ?
                             (7'h45) : (8'ha2)) < wire1) : ((&wire0) ^ wire1[(3'h6):(3'h5)])) : $signed(($signed((8'hbd)) ?
                         {wire2, wire4} : $signed(wire2)))) && (wire0 ?
                     $signed({$unsigned((8'h9f))}) : $signed(wire0[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      reg6 = $signed($signed((wire2[(5'h13):(5'h13)] == ($signed(wire3) ?
          $signed((8'hb4)) : (wire1 && wire0)))));
      for (forvar7 = (1'h0); (forvar7 < (2'h3)); forvar7 = (forvar7 + (1'h1)))
        begin
          if ($unsigned((8'had)))
            begin
              reg8 = reg6;
            end
          else
            begin
              reg9 <= (8'h9f);
              reg10 <= reg9[(1'h0):(1'h0)];
            end
          reg11 = $signed({$unsigned(reg6)});
        end
      if ($signed(wire0[(1'h1):(1'h0)]))
        begin
          if (reg9[(2'h2):(1'h0)])
            begin
              reg12 = ((8'haf) ? wire4[(4'h9):(3'h7)] : $unsigned(wire3));
            end
          else
            begin
              reg13 <= $signed((!reg9[(2'h2):(1'h0)]));
            end
          reg14 <= $unsigned({wire2});
          if (wire0)
            begin
              reg15 = ({(^~$unsigned(reg11))} ?
                  (!forvar7[(1'h0):(1'h0)]) : $signed({(reg8 || reg11[(2'h2):(1'h1)]),
                      $unsigned((~reg13))}));
              reg16 <= $signed(wire3[(4'hf):(4'h9)]);
            end
          else
            begin
              reg15 = (8'h9d);
              reg17 = $signed($signed((~(~|reg16))));
              reg18 <= (($unsigned($signed($signed(wire0))) && reg17) ?
                  (+(reg9[(1'h1):(1'h1)] + ($unsigned(reg11) ?
                      reg17[(4'h9):(4'h9)] : reg9[(2'h3):(2'h2)]))) : {wire0[(2'h3):(1'h0)]});
              reg19 = $unsigned(((&reg17[(1'h0):(1'h0)]) >= $unsigned(((!(8'h9d)) >>> $signed(reg13)))));
            end
          reg20 <= ((~&$unsigned(reg17)) ? wire4 : (-wire0));
        end
      else
        begin
          for (forvar12 = (1'h0); (forvar12 < (2'h3)); forvar12 = (forvar12 + (1'h1)))
            begin
              reg13 <= (reg9[(1'h1):(1'h0)] ?
                  $unsigned(($signed(((8'hbd) ?
                      reg11 : reg17)) + ((reg20 >= (8'hbe)) ?
                      wire1 : (forvar7 ? wire5 : reg18)))) : reg18);
              reg14 <= $unsigned(forvar12[(2'h2):(1'h0)]);
            end
          if (((^~reg18) ? reg20[(4'h9):(4'h8)] : $signed(wire3)))
            begin
              reg15 = {{$signed(wire0)}};
              reg17 = reg13[(4'ha):(4'h8)];
            end
          else
            begin
              reg16 <= {wire0[(3'h4):(1'h0)], reg16};
              reg18 <= (wire1[(3'h6):(1'h1)] ?
                  (reg20 && $unsigned(reg9)) : reg19);
              reg20 <= $signed(reg12);
              reg21 = {wire0};
            end
          for (forvar22 = (1'h0); (forvar22 < (3'h4)); forvar22 = (forvar22 + (1'h1)))
            begin
              reg23 = $signed((reg6[(2'h3):(2'h3)] ?
                  $unsigned(((~&wire0) ?
                      (wire2 ? (7'h48) : (7'h40)) : $signed(reg18))) : wire5));
              reg24 <= $unsigned((!$unsigned($unsigned((~^reg8)))));
            end
          reg25 <= {reg12, $unsigned($signed(((reg17 <= reg16) - (|reg13))))};
        end
      for (forvar26 = (1'h0); (forvar26 < (3'h4)); forvar26 = (forvar26 + (1'h1)))
        begin
          if (reg18)
            begin
              reg27 <= (^$signed(((&(reg10 >= reg20)) ~^ (~^$unsigned(reg21)))));
              reg28 = reg23[(1'h0):(1'h0)];
            end
          else
            begin
              reg27 <= (((|reg27[(1'h1):(1'h0)]) ?
                  (&{$signed((8'hb9)), (forvar7 & wire1)}) : (reg12 ?
                      $unsigned((~&reg18)) : ($unsigned(reg19) ?
                          (^~forvar12) : (reg28 && reg9)))) < (({reg8[(3'h5):(2'h3)]} ?
                  ((^reg13) && reg28[(1'h1):(1'h0)]) : (~$unsigned(reg12))) >= wire2));
              reg29 <= (^~$unsigned(($signed($unsigned(reg12)) ~^ (&(~|wire0)))));
              reg30 <= {(~|reg9[(2'h3):(2'h2)])};
            end
          reg31 <= reg13[(4'he):(4'h8)];
          reg32 = wire4[(2'h3):(1'h0)];
        end
    end
  assign wire33 = $signed({reg9[(3'h4):(2'h2)], (8'ha9)});
  assign wire34 = $signed(wire1[(1'h1):(1'h0)]);
  assign wire35 = (8'h9c);
  module36 #() modinst309 (.wire41(reg9), .wire37(reg10), .wire38(reg29), .wire39(reg24), .clk(clk), .wire40(wire4), .y(wire308));
  assign wire310 = reg24[(3'h6):(1'h1)];
  always
    @(posedge clk) begin
      reg311 <= (wire0[(2'h2):(2'h2)] && wire34);
      if ((~|wire4))
        begin
          for (forvar312 = (1'h0); (forvar312 < (2'h3)); forvar312 = (forvar312 + (1'h1)))
            begin
              reg313 = $unsigned({(|($unsigned(wire2) >> reg25[(5'h12):(4'hb)])),
                  $unsigned(((reg31 <= forvar312) > (reg30 >> (8'haa))))});
            end
          reg314 = (+((8'ha0) ? reg27[(2'h2):(1'h1)] : reg13));
        end
      else
        begin
          if ($unsigned((reg18[(4'h8):(3'h6)] ? (+reg18) : (~&reg13))))
            begin
              reg312 <= reg10[(1'h0):(1'h0)];
              reg313 = $unsigned((((8'hbf) || (|{reg18,
                  wire5})) < {$unsigned(reg18[(1'h1):(1'h1)]),
                  ((|wire0) >> $signed(wire1))}));
              reg315 <= (8'hac);
              reg316 <= $unsigned($signed((^~wire34[(4'h8):(4'h8)])));
              reg317 = (reg18 >= (((reg25[(1'h1):(1'h1)] > ((8'haf) ?
                      wire4 : reg311)) ?
                  ($signed((8'hbf)) ?
                      $signed(reg311) : wire0) : $unsigned((~|reg29))) * ((((8'ha2) != wire4) ?
                      $signed(reg313) : {reg13, reg315}) ?
                  (~&$signed(wire0)) : reg10)));
            end
          else
            begin
              reg313 = $unsigned((~(!((~reg316) ?
                  $unsigned((8'hb6)) : reg314))));
              reg315 <= (^~reg314[(4'hf):(2'h3)]);
              reg317 = (~|$signed(($unsigned(wire4[(4'hf):(4'hd)]) << wire5[(3'h6):(1'h1)])));
              reg318 <= (($signed(reg311) ?
                      (~|(~(reg24 >>> reg18))) : wire1[(4'ha):(4'ha)]) ?
                  (+reg312) : ({wire308[(1'h0):(1'h0)],
                      wire0[(1'h0):(1'h0)]} * ((~^(~wire5)) || ((!wire0) ?
                      reg27[(2'h2):(1'h1)] : (wire35 ? reg317 : wire2)))));
            end
          reg319 <= $unsigned($unsigned($unsigned((8'hb0))));
        end
      for (forvar320 = (1'h0); (forvar320 < (1'h0)); forvar320 = (forvar320 + (1'h1)))
        begin
          for (forvar321 = (1'h0); (forvar321 < (2'h2)); forvar321 = (forvar321 + (1'h1)))
            begin
              reg322 <= ((wire5 ? $signed((-(&reg315))) : $unsigned((8'ha7))) ?
                  $unsigned(reg313[(4'h8):(3'h6)]) : reg16[(5'h12):(2'h3)]);
              reg323 = $signed(wire2[(3'h6):(1'h1)]);
              reg324 = ({($unsigned((reg314 ?
                          reg27 : reg27)) <<< ($signed(wire34) < $signed(reg18)))} ?
                  ((8'hbc) ?
                      $signed($signed((8'hab))) : (8'hbc)) : ($unsigned($unsigned(((8'hba) + reg323))) | $signed({(reg319 && (8'ha5)),
                      reg27[(1'h0):(1'h0)]})));
              reg325 = (reg314 ?
                  ({(~|forvar312[(4'ha):(4'h9)]),
                      wire5[(4'h8):(3'h5)]} - ($signed((8'hb5)) || ($signed(wire33) ?
                      (8'hab) : (&wire34)))) : $unsigned($unsigned((~|(^~wire33)))));
            end
          for (forvar326 = (1'h0); (forvar326 < (2'h3)); forvar326 = (forvar326 + (1'h1)))
            begin
              reg327 = {wire5, wire308};
              reg328 <= reg323;
              reg329 <= $unsigned((reg27 != (&({forvar312, reg324} ?
                  $signed(wire2) : $signed(reg322)))));
              reg330 <= ($unsigned($unsigned(reg24)) ? forvar321 : wire5);
            end
        end
      if (reg313[(3'h7):(1'h0)])
        begin
          reg331 <= $signed((wire3[(4'hb):(1'h0)] ?
              (($unsigned(wire1) >= reg313[(3'h5):(3'h5)]) ?
                  (reg9[(3'h4):(1'h1)] ?
                      $signed(reg20) : (~&reg18)) : (wire0[(3'h4):(1'h1)] | (forvar321 ?
                      reg325 : reg324))) : $unsigned($signed((~^reg14)))));
          reg332 = (~(((&(wire308 >= reg24)) >> wire308[(3'h5):(2'h3)]) ?
              (8'ha7) : (wire1[(4'h8):(3'h7)] >> (reg10 ?
                  (~^reg27) : wire2[(4'hd):(4'h8)]))));
        end
      else
        begin
          for (forvar331 = (1'h0); (forvar331 < (3'h4)); forvar331 = (forvar331 + (1'h1)))
            begin
              reg333 <= $signed(reg328[(3'h6):(3'h6)]);
              reg334 = $signed(wire5[(5'h10):(4'h9)]);
              reg335 <= {reg315[(1'h1):(1'h0)]};
              reg336 = (8'ha5);
              reg337 <= ($unsigned(wire35) | (($unsigned((wire5 < reg323)) ?
                      reg315 : ((forvar312 != reg16) * ((8'ha5) || reg318))) ?
                  (!reg20[(1'h0):(1'h0)]) : ($signed((|reg29)) ?
                      reg336[(1'h0):(1'h0)] : $signed((~^reg318)))));
            end
          if ((~&$signed(reg327[(3'h5):(2'h3)])))
            begin
              reg338 = (7'h42);
              reg339 <= reg322;
            end
          else
            begin
              reg339 <= ({(~wire1[(1'h0):(1'h0)])} <<< (|(reg24[(4'h8):(3'h6)] ?
                  ($unsigned(wire1) ?
                      (reg314 ? wire3 : wire0) : reg315) : {reg14, reg335})));
              reg340 = $unsigned((reg316[(5'h12):(4'hc)] ?
                  ($signed((reg319 ?
                      wire35 : reg311)) ^ wire34[(4'ha):(3'h6)]) : (^$unsigned(wire3[(3'h7):(1'h0)]))));
            end
          if ($signed(($signed((^reg9)) <= (^$unsigned((&reg9))))))
            begin
              reg341 = $unsigned((^~$unsigned(reg333)));
              reg342 <= (forvar312 ~^ ((-({reg13, reg324} ?
                  $unsigned((7'h46)) : (wire35 ?
                      reg329 : forvar312))) + reg314[(3'h7):(2'h2)]));
            end
          else
            begin
              reg342 <= (~^(^~(wire310 >> $unsigned(reg341))));
              reg343 <= (!reg27[(2'h2):(1'h0)]);
              reg344 = wire4[(2'h2):(1'h0)];
              reg345 <= reg31;
              reg346 <= forvar320[(5'h11):(5'h10)];
            end
          if (reg340)
            begin
              reg347 <= wire1;
              reg348 <= $signed((reg334[(2'h3):(2'h2)] ^~ $signed($unsigned($signed(wire5)))));
              reg349 = (((reg325 ? {reg346, (^reg338)} : (~$unsigned(reg332))) ?
                  (^reg342[(1'h1):(1'h1)]) : (8'h9e)) - ({$unsigned(reg25)} ?
                  (((^~(8'hab)) ? forvar331[(2'h2):(1'h1)] : reg334) ?
                      reg345[(1'h1):(1'h1)] : {$unsigned(reg336),
                          $signed((7'h49))}) : $signed(reg27[(1'h0):(1'h0)])));
              reg350 <= forvar321;
              reg351 <= ($signed(wire34) == $unsigned(((8'haf) ^ ($signed(reg322) ?
                  reg328[(2'h2):(1'h0)] : $signed(reg328)))));
            end
          else
            begin
              reg347 <= reg345[(4'h9):(4'h8)];
              reg348 <= wire2;
            end
          reg352 = (~&($signed((!{reg324, reg16})) ?
              reg324[(1'h1):(1'h1)] : $unsigned($unsigned($unsigned((7'h40))))));
        end
    end
  module353 #() modinst469 (wire468, clk, reg20, reg16, reg14, reg331, reg31);
  assign wire470 = (reg25[(3'h4):(2'h3)] ?
                       ({wire1[(4'h8):(4'h8)]} || (reg10 ?
                           ($unsigned(reg9) ~^ $signed(reg329)) : ((~reg24) | $signed(reg29)))) : (~$signed($unsigned($signed((8'ha5))))));
  always
    @(posedge clk) begin
      reg471 <= (!(^wire468[(1'h1):(1'h0)]));
      reg472 = reg318[(2'h3):(2'h2)];
      reg473 = {(^~wire5),
          ((+((wire34 ? reg315 : reg330) < (!wire308))) ?
              reg20 : ((&$unsigned(reg319)) != $unsigned((reg31 ?
                  (8'ha0) : reg345))))};
      if ($unsigned((reg14[(4'hf):(4'hf)] ? (~^$signed((&reg333))) : (8'hb8))))
        begin
          reg474 <= $signed($signed((((reg322 | wire5) & $unsigned(wire0)) ?
              reg318[(1'h1):(1'h1)] : reg331)));
          reg475 <= $unsigned(reg31);
        end
      else
        begin
          reg474 <= (($signed((!$signed(reg16))) & wire5[(4'h9):(3'h4)]) <= $unsigned($signed($unsigned((reg31 & reg474)))));
        end
    end
  module476 #() modinst971 (wire970, clk, reg316, reg351, reg30, reg29, reg312);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module476
#(parameter param969 = (~|(~(~&(&((8'had) <= (8'ha2)))))))
(y, clk, wire481, wire480, wire479, wire478, wire477);
  output wire [(32'h47e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire481;
  input wire [(4'hf):(1'h0)] wire480;
  input wire signed [(4'h9):(1'h0)] wire479;
  input wire signed [(3'h4):(1'h0)] wire478;
  input wire signed [(4'ha):(1'h0)] wire477;
  wire signed [(3'h7):(1'h0)] wire915;
  wire [(5'h15):(1'h0)] wire532;
  wire [(3'h7):(1'h0)] wire530;
  wire signed [(5'h12):(1'h0)] wire506;
  wire [(4'hd):(1'h0)] wire482;
  wire signed [(5'h16):(1'h0)] wire917;
  wire [(4'hf):(1'h0)] wire918;
  wire signed [(2'h3):(1'h0)] wire919;
  wire signed [(4'ha):(1'h0)] wire920;
  wire signed [(4'h8):(1'h0)] wire921;
  wire [(5'h15):(1'h0)] wire965;
  reg [(5'h10):(1'h0)] reg968 = (1'h0);
  reg [(4'ha):(1'h0)] reg531 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg529 = (1'h0);
  reg [(3'h4):(1'h0)] reg528 = (1'h0);
  reg [(4'h9):(1'h0)] reg526 = (1'h0);
  reg [(5'h10):(1'h0)] reg522 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg521 = (1'h0);
  reg [(5'h18):(1'h0)] reg520 = (1'h0);
  reg [(5'h10):(1'h0)] reg519 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg517 = (1'h0);
  reg [(5'h11):(1'h0)] reg516 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg515 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg512 = (1'h0);
  reg [(4'ha):(1'h0)] reg511 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg509 = (1'h0);
  reg [(4'ha):(1'h0)] reg505 = (1'h0);
  reg [(5'h16):(1'h0)] reg504 = (1'h0);
  reg [(5'h18):(1'h0)] reg500 = (1'h0);
  reg [(4'hd):(1'h0)] reg499 = (1'h0);
  reg [(4'hf):(1'h0)] reg497 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg494 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg493 = (1'h0);
  reg [(5'h13):(1'h0)] reg491 = (1'h0);
  reg [(4'h9):(1'h0)] reg490 = (1'h0);
  reg [(5'h16):(1'h0)] reg489 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg487 = (1'h0);
  reg [(4'hb):(1'h0)] reg485 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg484 = (1'h0);
  reg [(3'h6):(1'h0)] reg483 = (1'h0);
  reg [(3'h4):(1'h0)] reg923 = (1'h0);
  reg [(4'hd):(1'h0)] reg928 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg929 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg934 = (1'h0);
  reg [(5'h18):(1'h0)] reg936 = (1'h0);
  reg [(4'h9):(1'h0)] reg941 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg943 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg944 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg946 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg967 = (1'h0);
  reg signed [(4'he):(1'h0)] reg945 = (1'h0);
  reg [(5'h17):(1'h0)] reg942 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg940 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar939 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg938 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg937 = (1'h0);
  reg [(4'hd):(1'h0)] forvar935 = (1'h0);
  reg [(4'h9):(1'h0)] reg933 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg932 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar931 = (1'h0);
  reg [(5'h18):(1'h0)] forvar930 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg927 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg926 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg925 = (1'h0);
  reg [(5'h13):(1'h0)] reg924 = (1'h0);
  reg [(5'h17):(1'h0)] reg922 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg527 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar525 = (1'h0);
  reg [(4'hf):(1'h0)] reg524 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar523 = (1'h0);
  reg signed [(4'he):(1'h0)] reg518 = (1'h0);
  reg [(2'h2):(1'h0)] forvar514 = (1'h0);
  reg [(2'h2):(1'h0)] reg513 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg510 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg508 = (1'h0);
  reg [(3'h6):(1'h0)] forvar507 = (1'h0);
  reg [(5'h11):(1'h0)] reg503 = (1'h0);
  reg [(2'h3):(1'h0)] reg502 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg501 = (1'h0);
  reg [(4'hb):(1'h0)] reg498 = (1'h0);
  reg [(5'h15):(1'h0)] forvar483 = (1'h0);
  reg [(5'h12):(1'h0)] reg496 = (1'h0);
  reg [(5'h11):(1'h0)] reg495 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg492 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg488 = (1'h0);
  reg [(3'h6):(1'h0)] reg486 = (1'h0);
  assign y = {wire915,
                 wire532,
                 wire530,
                 wire506,
                 wire482,
                 wire917,
                 wire918,
                 wire919,
                 wire920,
                 wire921,
                 wire965,
                 reg968,
                 reg531,
                 reg529,
                 reg528,
                 reg526,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg517,
                 reg516,
                 reg515,
                 reg512,
                 reg511,
                 reg509,
                 reg505,
                 reg504,
                 reg500,
                 reg499,
                 reg497,
                 reg494,
                 reg493,
                 reg491,
                 reg490,
                 reg489,
                 reg487,
                 reg485,
                 reg484,
                 reg483,
                 reg923,
                 reg928,
                 reg929,
                 reg934,
                 reg936,
                 reg941,
                 reg943,
                 reg944,
                 reg946,
                 reg967,
                 reg945,
                 reg942,
                 reg940,
                 forvar939,
                 reg938,
                 reg937,
                 forvar935,
                 reg933,
                 reg932,
                 forvar931,
                 forvar930,
                 reg927,
                 reg926,
                 reg925,
                 reg924,
                 reg922,
                 reg527,
                 forvar525,
                 reg524,
                 forvar523,
                 reg518,
                 forvar514,
                 reg513,
                 reg510,
                 reg508,
                 forvar507,
                 reg503,
                 reg502,
                 reg501,
                 reg498,
                 forvar483,
                 reg496,
                 reg495,
                 reg492,
                 reg488,
                 reg486,
                 (1'h0)};
  assign wire482 = (~&(~(wire480 + $signed(wire477))));
  always
    @(posedge clk) begin
      if ($signed($unsigned(wire477)))
        begin
          reg483 <= $unsigned((~$unsigned($signed($signed(wire480)))));
          if (((wire480 >>> ({(|wire477),
              (wire477 ?
                  wire478 : (7'h49))} & $unsigned(wire478))) > wire482[(1'h1):(1'h1)]))
            begin
              reg484 <= (8'hb2);
              reg485 <= $unsigned((!(~^(8'ha3))));
            end
          else
            begin
              reg486 = ({(-wire481),
                  ($signed(wire482[(1'h0):(1'h0)]) != {$unsigned(wire477),
                      wire478})} != ($unsigned($unsigned($signed(reg483))) ?
                  $signed(reg483[(1'h1):(1'h1)]) : wire477));
              reg487 <= ((+((-(7'h45)) ?
                      {(~^wire480)} : ((wire478 >>> wire479) >= (!wire482)))) ?
                  (-((!(~reg485)) ^ wire480)) : ((+$signed($signed(reg486))) < ({(~wire480)} ?
                      (-(wire480 - wire479)) : (^~wire482))));
              reg488 = reg484;
              reg489 <= ((^~(!$signed($signed(reg485)))) * {((~^(wire480 != reg483)) >> {$signed(wire482)})});
            end
          if (wire478[(1'h1):(1'h0)])
            begin
              reg490 <= ($signed(((~&reg486[(3'h6):(1'h1)]) ~^ $unsigned(((8'hb7) ?
                      wire481 : reg484)))) ?
                  $signed(reg485) : {$unsigned(wire480[(2'h3):(2'h2)])});
              reg491 <= (((~&$signed({wire478,
                      (8'hae)})) * reg485[(3'h7):(3'h6)]) ?
                  {((~^$signed(reg487)) ?
                          (((8'hb1) == reg488) ?
                              $signed(reg483) : reg488[(3'h6):(3'h5)]) : ((&reg485) ?
                              $signed((8'ha0)) : {reg487,
                                  wire481}))} : ($unsigned(($signed(reg485) ?
                      wire480 : $signed(reg484))) << (($unsigned(reg488) ?
                          $signed(wire477) : $unsigned(reg488)) ?
                      wire482 : $unsigned(reg484[(4'hf):(4'he)]))));
              reg492 = reg484;
              reg493 <= (reg492[(2'h3):(2'h2)] >> $unsigned($unsigned({{reg483,
                      reg485}})));
              reg494 <= reg486[(3'h6):(1'h1)];
            end
          else
            begin
              reg492 = (($signed(wire480) <= $unsigned(({reg494} ?
                      wire478 : (~^reg493)))) ?
                  $signed($signed($signed((reg491 + wire480)))) : ({$unsigned((~|wire478)),
                      $signed((reg490 < wire481))} != wire477));
              reg495 = $signed((7'h49));
              reg496 = {(~|((wire482[(1'h0):(1'h0)] <= (reg495 < reg489)) ?
                      (-(reg485 ? (7'h48) : reg487)) : reg485)),
                  {$unsigned((!wire477[(2'h3):(2'h3)])), wire481}};
            end
        end
      else
        begin
          for (forvar483 = (1'h0); (forvar483 < (1'h1)); forvar483 = (forvar483 + (1'h1)))
            begin
              reg484 <= wire478[(2'h2):(2'h2)];
              reg485 <= {reg496[(5'h10):(4'he)]};
            end
        end
      if (wire482[(3'h5):(3'h5)])
        begin
          if (reg488[(1'h1):(1'h0)])
            begin
              reg497 <= ($signed((($signed((8'hb7)) == $unsigned(reg485)) == reg496)) ?
                  $unsigned($signed($signed((wire481 != wire478)))) : ((|$unsigned((reg486 ?
                          reg491 : (7'h40)))) ?
                      (7'h40) : $signed($signed(reg494[(1'h0):(1'h0)]))));
              reg498 = (($unsigned(((+reg491) ? (^(8'ha5)) : (8'hbf))) ?
                      wire481 : {reg494}) ?
                  wire482[(1'h0):(1'h0)] : (|(~reg487[(4'ha):(4'h9)])));
              reg499 <= reg497;
              reg500 <= $unsigned((((^{reg490}) ?
                  ((reg493 & wire481) | wire477) : $unsigned((reg492 ?
                      reg498 : reg496))) <<< $signed(((!reg496) <= $unsigned(reg489)))));
            end
          else
            begin
              reg498 = ($unsigned((^~$signed((wire477 + wire478)))) ?
                  {(((reg485 <<< reg499) == reg487[(4'h8):(3'h4)]) < reg493[(4'h8):(1'h0)])} : $signed({$signed((reg494 >> (8'hb6)))}));
              reg501 = (!($signed((reg486[(2'h2):(2'h2)] ?
                  reg499[(2'h3):(2'h2)] : {reg490,
                      (8'ha7)})) || {wire479[(3'h6):(3'h6)],
                  ($signed(reg499) ^~ (reg491 >>> wire482))}));
              reg502 = $unsigned(reg496);
              reg503 = (8'hba);
              reg504 <= reg493;
            end
        end
      else
        begin
          reg497 <= ($unsigned(reg497[(3'h5):(3'h5)]) != wire478);
          reg499 <= {$signed(((~^((8'hb2) ? reg483 : (7'h45))) < reg494)),
              $unsigned((reg486[(3'h5):(3'h5)] ?
                  reg500 : reg501[(2'h3):(1'h1)]))};
          reg500 <= ($unsigned($unsigned($unsigned(((8'hae) ?
              reg493 : reg502)))) && ((reg494 ?
              reg492 : {(!reg485)}) ^ $unsigned(reg501[(2'h3):(1'h0)])));
        end
      reg505 <= (-(~^$signed((~$signed((8'ha5))))));
    end
  assign wire506 = $signed(reg499[(4'h8):(3'h7)]);
  always
    @(posedge clk) begin
      for (forvar507 = (1'h0); (forvar507 < (2'h3)); forvar507 = (forvar507 + (1'h1)))
        begin
          if ($signed(reg487))
            begin
              reg508 = $unsigned((reg491[(2'h2):(1'h0)] ~^ {$signed(forvar507),
                  reg489}));
              reg509 <= reg494[(3'h6):(3'h6)];
            end
          else
            begin
              reg508 = (+$signed(reg494));
              reg510 = ((reg500 - (((reg504 ? (8'hb5) : wire482) ?
                          reg485 : reg504) ?
                      ($unsigned((8'ha2)) ^ (reg483 == reg484)) : (wire480[(3'h4):(2'h3)] >> $signed(wire478)))) ?
                  reg508 : (wire506[(5'h11):(1'h0)] <<< reg497));
              reg511 <= $signed((~|$signed(({reg505, wire506} ?
                  reg499 : (reg509 ? wire479 : wire481)))));
              reg512 <= reg491[(2'h3):(2'h3)];
              reg513 = (reg497 ?
                  reg484[(3'h7):(1'h1)] : (-($signed($unsigned(reg500)) ?
                      $signed($unsigned((7'h40))) : ($signed(reg499) ?
                          $unsigned(reg505) : $signed(reg485)))));
            end
          for (forvar514 = (1'h0); (forvar514 < (1'h0)); forvar514 = (forvar514 + (1'h1)))
            begin
              reg515 <= wire480;
              reg516 <= $signed($signed((^~((-(8'hbc)) - $signed(wire478)))));
              reg517 <= (^reg510);
            end
          if ($unsigned((reg504 >= $signed(($signed(reg493) ?
              (wire480 ? reg483 : (8'ha5)) : reg516[(4'he):(1'h1)])))))
            begin
              reg518 = ((|($signed((reg516 | (8'hbe))) ^ ($unsigned(forvar507) ?
                      (^wire481) : (reg483 - (8'h9f))))) ?
                  reg513[(2'h2):(1'h0)] : (~^(|$signed(wire482[(3'h5):(3'h5)]))));
              reg519 <= $unsigned({{$unsigned((wire480 - (7'h40))),
                      ($signed(reg489) | (&reg490))}});
            end
          else
            begin
              reg519 <= (&(^~((((8'hbd) ?
                  reg518 : reg497) != (reg490 < wire479)) - ((reg485 * reg490) | (-(8'h9e))))));
              reg520 <= (~|(reg490[(3'h7):(2'h2)] ?
                  $unsigned($unsigned((reg493 ?
                      (8'hb9) : wire478))) : reg484[(4'hb):(2'h3)]));
              reg521 <= forvar507[(1'h1):(1'h1)];
              reg522 <= $unsigned(((((reg499 ^ reg504) & (8'ha8)) ?
                  ((wire480 + reg515) | (+reg483)) : (~(reg487 ?
                      reg512 : reg500))) <<< $unsigned(reg483)));
            end
          for (forvar523 = (1'h0); (forvar523 < (2'h3)); forvar523 = (forvar523 + (1'h1)))
            begin
              reg524 = reg499;
            end
          for (forvar525 = (1'h0); (forvar525 < (2'h3)); forvar525 = (forvar525 + (1'h1)))
            begin
              reg526 <= (((^$unsigned((reg491 ?
                      (8'ha4) : forvar523))) >= reg518[(2'h2):(1'h1)]) ?
                  $unsigned(wire482) : (reg483 && $signed($unsigned(reg512))));
              reg527 = {$signed(reg485), $unsigned((^~reg516))};
            end
        end
      reg528 <= (($signed((reg516[(3'h7):(2'h3)] ?
              reg499[(4'hb):(4'ha)] : {reg509})) ?
          reg499 : reg511[(1'h1):(1'h1)]) > reg516[(2'h2):(1'h0)]);
      reg529 <= $signed($unsigned((+(reg515 ?
          ((7'h40) >= reg511) : $unsigned((8'hbe))))));
    end
  assign wire530 = $unsigned((~&(($signed(wire480) ^~ (-reg493)) ?
                       (&$unsigned(reg517)) : $signed((reg489 ?
                           (8'had) : reg515)))));
  always
    @(posedge clk) begin
      reg531 <= $unsigned(reg487);
    end
  assign wire532 = (~|{($signed($unsigned(reg516)) & $unsigned(reg483[(1'h1):(1'h0)])),
                       ((|(reg512 ? reg522 : reg499)) ^ reg511)});
  module533 #() modinst916 (.y(wire915), .wire537(reg485), .wire534(reg484), .wire536(reg515), .clk(clk), .wire535(wire482));
  assign wire917 = ({$signed({$unsigned((8'had)), $signed(reg484)}),
                           ($signed($signed(reg517)) ^~ $unsigned($signed(reg516)))} ?
                       ($unsigned(reg497) ~^ $signed($unsigned((~^(7'h49))))) : ($unsigned($unsigned({reg499})) ?
                           $signed($unsigned(((8'hbc) ?
                               wire506 : reg497))) : ($unsigned($unsigned(wire482)) ?
                               wire532[(5'h15):(4'ha)] : {$unsigned(wire480),
                                   $signed(reg522)})));
  assign wire918 = reg517;
  assign wire919 = {(~((reg487[(4'ha):(2'h3)] - {wire918}) ?
                           ((8'hb5) ?
                               $unsigned(reg522) : wire477[(4'h9):(4'h8)]) : wire481))};
  assign wire920 = wire530;
  assign wire921 = reg519;
  always
    @(posedge clk) begin
      reg922 = (~&reg505[(4'ha):(1'h1)]);
      if (reg515)
        begin
          reg923 <= $unsigned(($signed($signed((8'ha8))) * $unsigned(($signed(wire919) ?
              {reg529, reg493} : (wire478 ? reg484 : reg493)))));
        end
      else
        begin
          reg924 = $unsigned(reg494);
          reg925 = (^~reg511[(2'h2):(2'h2)]);
          reg926 = (~&({((reg517 ? (8'hb4) : reg528) & (wire481 ?
                  reg512 : wire506)),
              ((^reg529) - $signed(reg500))} ~^ {(&((8'hbf) ? reg515 : reg924)),
              reg521[(5'h18):(4'hd)]}));
          reg927 = (8'hbf);
        end
      reg928 <= (|(-reg504[(2'h3):(2'h2)]));
      reg929 <= $unsigned(((((~|reg483) != (^reg511)) ?
              $signed(reg489[(5'h11):(4'ha)]) : $unsigned((reg497 ?
                  (8'hb4) : reg500))) ?
          $signed(($unsigned((8'hac)) ?
              $signed((8'hb1)) : {reg490})) : {wire530[(3'h4):(3'h4)],
              $unsigned(wire482)}));
      for (forvar930 = (1'h0); (forvar930 < (3'h4)); forvar930 = (forvar930 + (1'h1)))
        begin
          for (forvar931 = (1'h0); (forvar931 < (1'h1)); forvar931 = (forvar931 + (1'h1)))
            begin
              reg932 = ($signed(($signed((+reg924)) >> (((8'hbf) ?
                      wire478 : reg500) <= (8'hbf)))) ?
                  (forvar931 ?
                      ((+reg491[(3'h5):(2'h3)]) ^ reg929) : $unsigned((~^(wire480 <<< reg511)))) : reg924[(2'h3):(2'h3)]);
              reg933 = wire479;
              reg934 <= (|(^($signed($unsigned(wire920)) ?
                  (reg528[(2'h3):(2'h3)] ?
                      (^~reg512) : $unsigned(reg515)) : (|$unsigned(reg505)))));
            end
          for (forvar935 = (1'h0); (forvar935 < (3'h4)); forvar935 = (forvar935 + (1'h1)))
            begin
              reg936 <= (reg493[(3'h6):(3'h5)] || ({$signed((7'h47))} ?
                  $signed($signed((+wire920))) : $unsigned((~&$unsigned((7'h45))))));
              reg937 = reg928;
              reg938 = (7'h44);
            end
          for (forvar939 = (1'h0); (forvar939 < (3'h4)); forvar939 = (forvar939 + (1'h1)))
            begin
              reg940 = ((($signed((reg489 >> wire506)) ?
                      $signed(reg923) : ((!reg512) & reg520)) ?
                  (|((+wire530) >> $unsigned((8'hb7)))) : (7'h46)) || ($signed((~&$signed(reg924))) ?
                  (((forvar930 ? reg519 : wire917) ? (7'h49) : reg512) ?
                      wire921[(1'h1):(1'h0)] : reg511) : (8'hb3)));
              reg941 <= {forvar930, wire915};
              reg942 = (^~(~&reg932[(5'h15):(5'h13)]));
              reg943 <= {(-(wire915[(2'h3):(2'h3)] ?
                      wire918[(4'h8):(1'h1)] : (8'hab)))};
              reg944 <= wire917;
            end
          reg945 = ({(|{(8'haf), reg485})} ? reg512 : $unsigned(reg933));
          reg946 <= ($signed((((+reg520) ?
                      $signed(wire919) : (wire479 < wire915)) ?
                  wire915[(1'h1):(1'h1)] : {$signed(reg928)})) ?
              {$signed((^{reg928, reg927})),
                  $signed($signed(reg922))} : wire530[(2'h3):(2'h2)]);
        end
    end
  module947 #() modinst966 (.clk(clk), .y(wire965), .wire948(reg944), .wire951(reg493), .wire950(wire480), .wire949(reg489));
  always
    @(posedge clk) begin
      reg967 = reg485;
      reg968 <= $unsigned(({reg509} == ((8'haa) >= $signed((wire915 ?
          reg509 : reg944)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module353
#(parameter param466 = ((&(~((8'hae) ? ((8'h9e) ? (7'h48) : (7'h44)) : {(8'ha3)}))) <= ({((~(8'ha1)) << ((7'h40) << (8'h9e))), (~|(^(8'h9f)))} - ((~&((8'ha0) ? (7'h46) : (8'hb3))) ? {((7'h46) + (8'hbc))} : {((8'ha6) ? (8'hb9) : (7'h41)), (~(8'hbb))}))), 
parameter param467 = ((~&{(~&(param466 | param466)), (|{param466, param466})}) ? (-param466) : (8'ha5)))
(y, clk, wire358, wire357, wire356, wire355, wire354);
  output wire [(32'h5a9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h7):(1'h0)] wire358;
  input wire signed [(2'h2):(1'h0)] wire357;
  input wire [(4'hf):(1'h0)] wire356;
  input wire signed [(2'h2):(1'h0)] wire355;
  input wire [(2'h3):(1'h0)] wire354;
  wire signed [(5'h13):(1'h0)] wire452;
  wire signed [(5'h14):(1'h0)] wire451;
  wire signed [(5'h17):(1'h0)] wire377;
  reg [(3'h6):(1'h0)] reg465 = (1'h0);
  reg [(4'h9):(1'h0)] reg464 = (1'h0);
  reg [(5'h11):(1'h0)] reg462 = (1'h0);
  reg [(5'h10):(1'h0)] reg460 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg457 = (1'h0);
  reg [(5'h13):(1'h0)] reg449 = (1'h0);
  reg [(5'h17):(1'h0)] reg446 = (1'h0);
  reg [(2'h3):(1'h0)] reg443 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg442 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg440 = (1'h0);
  reg [(4'h8):(1'h0)] reg435 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg433 = (1'h0);
  reg [(5'h11):(1'h0)] reg431 = (1'h0);
  reg [(2'h3):(1'h0)] reg430 = (1'h0);
  reg [(3'h6):(1'h0)] reg428 = (1'h0);
  reg [(4'he):(1'h0)] reg426 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg424 = (1'h0);
  reg [(2'h2):(1'h0)] reg423 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg421 = (1'h0);
  reg [(4'ha):(1'h0)] reg418 = (1'h0);
  reg [(5'h14):(1'h0)] reg417 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg412 = (1'h0);
  reg [(3'h4):(1'h0)] reg408 = (1'h0);
  reg [(4'h9):(1'h0)] reg407 = (1'h0);
  reg [(2'h2):(1'h0)] reg403 = (1'h0);
  reg [(4'hb):(1'h0)] reg402 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg401 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg398 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg396 = (1'h0);
  reg [(5'h10):(1'h0)] reg395 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg390 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg389 = (1'h0);
  reg [(2'h2):(1'h0)] reg387 = (1'h0);
  reg [(5'h11):(1'h0)] reg386 = (1'h0);
  reg [(4'ha):(1'h0)] reg384 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg381 = (1'h0);
  reg [(4'hf):(1'h0)] reg379 = (1'h0);
  reg [(4'hf):(1'h0)] reg370 = (1'h0);
  reg [(3'h4):(1'h0)] reg369 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg367 = (1'h0);
  reg [(4'hf):(1'h0)] reg364 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg361 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg360 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg463 = (1'h0);
  reg [(5'h10):(1'h0)] reg461 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg459 = (1'h0);
  reg [(3'h4):(1'h0)] forvar458 = (1'h0);
  reg [(4'hf):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar455 = (1'h0);
  reg [(2'h3):(1'h0)] reg454 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar453 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg450 = (1'h0);
  reg signed [(4'he):(1'h0)] reg448 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg447 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg445 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg444 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg441 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg439 = (1'h0);
  reg [(5'h10):(1'h0)] reg438 = (1'h0);
  reg [(5'h10):(1'h0)] reg437 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg436 = (1'h0);
  reg [(5'h10):(1'h0)] reg434 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg432 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg429 = (1'h0);
  reg [(4'hd):(1'h0)] reg427 = (1'h0);
  reg [(5'h17):(1'h0)] forvar425 = (1'h0);
  reg [(5'h18):(1'h0)] forvar422 = (1'h0);
  reg [(5'h15):(1'h0)] reg420 = (1'h0);
  reg [(2'h2):(1'h0)] forvar419 = (1'h0);
  reg [(4'h9):(1'h0)] reg415 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg414 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar413 = (1'h0);
  reg [(3'h4):(1'h0)] forvar411 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar410 = (1'h0);
  reg [(5'h15):(1'h0)] reg406 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar405 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg397 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg409 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar406 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg405 = (1'h0);
  reg [(4'hb):(1'h0)] reg404 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg400 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar399 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar397 = (1'h0);
  reg [(4'hc):(1'h0)] forvar391 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar387 = (1'h0);
  reg [(4'hc):(1'h0)] forvar384 = (1'h0);
  reg [(5'h11):(1'h0)] reg394 = (1'h0);
  reg [(4'hb):(1'h0)] reg393 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg392 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg391 = (1'h0);
  reg [(2'h3):(1'h0)] reg388 = (1'h0);
  reg [(2'h2):(1'h0)] reg385 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg383 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg382 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar380 = (1'h0);
  reg [(5'h10):(1'h0)] reg378 = (1'h0);
  reg [(4'he):(1'h0)] reg376 = (1'h0);
  reg [(4'hd):(1'h0)] reg375 = (1'h0);
  reg [(2'h2):(1'h0)] reg374 = (1'h0);
  reg [(5'h17):(1'h0)] forvar373 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg372 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar371 = (1'h0);
  reg [(5'h14):(1'h0)] reg368 = (1'h0);
  reg [(4'hf):(1'h0)] reg366 = (1'h0);
  reg [(4'ha):(1'h0)] reg365 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar362 = (1'h0);
  reg [(5'h15):(1'h0)] reg359 = (1'h0);
  assign y = {wire452,
                 wire451,
                 wire377,
                 reg465,
                 reg464,
                 reg462,
                 reg460,
                 reg457,
                 reg449,
                 reg446,
                 reg443,
                 reg442,
                 reg440,
                 reg435,
                 reg433,
                 reg431,
                 reg430,
                 reg428,
                 reg426,
                 reg424,
                 reg423,
                 reg421,
                 reg418,
                 reg417,
                 reg416,
                 reg412,
                 reg408,
                 reg407,
                 reg403,
                 reg402,
                 reg401,
                 reg398,
                 reg396,
                 reg395,
                 reg390,
                 reg389,
                 reg387,
                 reg386,
                 reg384,
                 reg381,
                 reg379,
                 reg370,
                 reg369,
                 reg367,
                 reg364,
                 reg361,
                 reg360,
                 reg463,
                 reg461,
                 reg459,
                 forvar458,
                 reg456,
                 forvar455,
                 reg454,
                 forvar453,
                 reg450,
                 reg448,
                 reg447,
                 reg445,
                 reg444,
                 reg441,
                 reg439,
                 reg438,
                 reg437,
                 reg436,
                 reg434,
                 reg432,
                 reg429,
                 reg427,
                 forvar425,
                 forvar422,
                 reg420,
                 forvar419,
                 reg415,
                 reg414,
                 forvar413,
                 forvar411,
                 forvar410,
                 reg406,
                 forvar405,
                 reg397,
                 reg409,
                 forvar406,
                 reg405,
                 reg404,
                 reg400,
                 forvar399,
                 forvar397,
                 forvar391,
                 forvar387,
                 forvar384,
                 reg394,
                 reg393,
                 reg392,
                 reg391,
                 reg388,
                 reg385,
                 reg383,
                 reg382,
                 forvar380,
                 reg378,
                 reg376,
                 reg375,
                 reg374,
                 forvar373,
                 reg372,
                 forvar371,
                 reg368,
                 reg366,
                 reg365,
                 reg363,
                 forvar362,
                 reg359,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg359 = ({(wire356[(4'h9):(3'h5)] ? wire355 : wire354[(2'h3):(2'h3)]),
          $signed((((8'hba) ?
              wire357 : wire355) ^~ $unsigned(wire354)))} <<< wire357[(2'h2):(2'h2)]);
      reg360 <= $unsigned((+(^((^wire357) ?
          $signed(wire358) : (wire354 ? wire356 : wire358)))));
    end
  always
    @(posedge clk) begin
      reg361 <= ((~^(wire357[(1'h0):(1'h0)] ?
              ($unsigned((8'hbb)) <= (~^reg360)) : {{wire355, wire356}})) ?
          wire357[(1'h0):(1'h0)] : (wire354 >>> $unsigned($unsigned({(7'h44)}))));
      for (forvar362 = (1'h0); (forvar362 < (2'h3)); forvar362 = (forvar362 + (1'h1)))
        begin
          reg363 = ($unsigned((!wire357)) != (~&forvar362[(1'h1):(1'h1)]));
          reg364 <= $unsigned(wire357[(2'h2):(1'h0)]);
          reg365 = reg363;
          reg366 = ((|reg361[(2'h3):(1'h0)]) - $signed($signed($unsigned((wire355 + reg364)))));
          reg367 <= $unsigned(((~|wire354) ?
              (|(~|$unsigned(wire358))) : ($signed((reg360 ?
                  reg361 : reg360)) == reg363[(3'h7):(3'h5)])));
        end
    end
  always
    @(posedge clk) begin
      reg368 = ((~((wire355[(2'h2):(2'h2)] ?
          $signed(wire355) : reg364[(3'h4):(1'h1)]) ^~ (8'hbc))) * reg367[(2'h3):(1'h1)]);
      reg369 <= $signed($unsigned($unsigned($signed((wire356 >= reg368)))));
      reg370 <= reg360;
    end
  always
    @(posedge clk) begin
      for (forvar371 = (1'h0); (forvar371 < (1'h0)); forvar371 = (forvar371 + (1'h1)))
        begin
          reg372 = {(~|$signed(reg369)), {wire355}};
          for (forvar373 = (1'h0); (forvar373 < (3'h4)); forvar373 = (forvar373 + (1'h1)))
            begin
              reg374 = (wire357[(2'h2):(2'h2)] ^~ $unsigned($unsigned($signed((^reg361)))));
            end
          reg375 = forvar371;
        end
      reg376 = wire354[(1'h0):(1'h0)];
    end
  assign wire377 = $unsigned(($unsigned(($unsigned((8'ha4)) ?
                           (~&reg369) : wire355)) ?
                       $signed(($signed(reg364) ?
                           (wire356 * wire356) : (^~reg367))) : ({$signed(reg370)} & reg364)));
  always
    @(posedge clk) begin
      reg378 = reg364[(1'h1):(1'h1)];
      reg379 <= wire355[(1'h0):(1'h0)];
      for (forvar380 = (1'h0); (forvar380 < (3'h4)); forvar380 = (forvar380 + (1'h1)))
        begin
          reg381 <= wire354[(1'h1):(1'h1)];
          reg382 = wire357[(1'h0):(1'h0)];
          reg383 = (|$signed((($signed((7'h49)) ?
              {wire355} : reg379[(4'hc):(4'ha)]) >= $unsigned((wire355 ?
              wire355 : wire356)))));
        end
      if ((forvar380[(1'h1):(1'h1)] - $unsigned(wire355)))
        begin
          if ((~|$signed($signed(($signed((8'h9c)) ?
              (!reg378) : (reg361 >= reg367))))))
            begin
              reg384 <= {wire377};
              reg385 = wire357[(1'h1):(1'h0)];
            end
          else
            begin
              reg384 <= $unsigned(($signed((&(wire358 ? reg381 : wire357))) ?
                  $unsigned((~^$unsigned(reg383))) : reg360[(1'h1):(1'h1)]));
              reg386 <= $signed(reg385[(1'h0):(1'h0)]);
              reg387 <= $signed(reg364);
              reg388 = (wire354[(2'h3):(1'h1)] >>> reg387[(1'h0):(1'h0)]);
              reg389 <= {((~|reg370) ~^ wire355), reg360};
            end
          if (reg384[(2'h2):(1'h1)])
            begin
              reg390 <= (((reg386 + ($unsigned(reg370) ? {(8'ha9)} : reg379)) ?
                  reg388 : $signed($signed((wire358 >> wire377)))) >= (^~(reg370[(3'h7):(1'h1)] + $signed((reg381 && reg386)))));
              reg391 = (7'h43);
            end
          else
            begin
              reg390 <= reg390;
              reg391 = reg382[(4'hb):(3'h7)];
              reg392 = {$signed((($signed(reg385) || reg361[(1'h0):(1'h0)]) > reg367)),
                  $unsigned(({reg369} > ((wire357 ?
                      reg386 : reg385) <<< (|reg367))))};
              reg393 = $signed($unsigned(({(reg370 ? reg390 : reg378)} ?
                  (!reg392[(5'h14):(1'h1)]) : $signed(reg387[(1'h1):(1'h0)]))));
              reg394 = $unsigned(reg392[(1'h1):(1'h0)]);
            end
        end
      else
        begin
          for (forvar384 = (1'h0); (forvar384 < (2'h3)); forvar384 = (forvar384 + (1'h1)))
            begin
              reg385 = reg361[(1'h1):(1'h1)];
            end
          reg386 <= {{reg394[(4'hf):(4'he)],
                  (((~(8'had)) && $signed(reg387)) <= reg381[(3'h5):(3'h4)])}};
          for (forvar387 = (1'h0); (forvar387 < (1'h1)); forvar387 = (forvar387 + (1'h1)))
            begin
              reg389 <= (reg379 ?
                  ({$unsigned((wire358 - (8'hb2))),
                          {((8'hac) * reg387), {reg382}}} ?
                      (-forvar384) : (^~wire354)) : reg360[(2'h2):(1'h0)]);
              reg390 <= reg361;
            end
          for (forvar391 = (1'h0); (forvar391 < (3'h4)); forvar391 = (forvar391 + (1'h1)))
            begin
              reg392 = (^~(~|{$unsigned(reg361[(1'h1):(1'h1)]),
                  {(reg389 ? reg387 : forvar387)}}));
            end
        end
    end
  always
    @(posedge clk) begin
      reg395 <= (((~wire357[(1'h0):(1'h0)]) ?
              (reg367[(3'h6):(2'h3)] <= $signed($signed(wire358))) : reg381[(4'h9):(4'h8)]) ?
          ((wire358 ? $signed($unsigned(reg390)) : reg384) ?
              (($unsigned(wire354) == reg384) * (reg390 ?
                  {(7'h40)} : (reg369 >> reg369))) : (~&($unsigned(wire377) != reg367[(3'h6):(2'h2)]))) : $unsigned((^((reg381 ?
              reg386 : (8'hb1)) >>> reg379[(4'hf):(2'h3)]))));
      if (reg384)
        begin
          reg396 <= reg379;
          for (forvar397 = (1'h0); (forvar397 < (3'h4)); forvar397 = (forvar397 + (1'h1)))
            begin
              reg398 <= (~((({(8'haa)} == $unsigned(reg367)) && ((wire356 ?
                      reg381 : reg379) ^ (~^forvar397))) ?
                  reg384[(4'h8):(1'h0)] : ($signed(reg361) ?
                      reg379[(4'hb):(3'h5)] : $unsigned($signed(reg395)))));
            end
          for (forvar399 = (1'h0); (forvar399 < (2'h3)); forvar399 = (forvar399 + (1'h1)))
            begin
              reg400 = reg364[(4'he):(3'h4)];
              reg401 <= (^((({(8'haa), (8'hb6)} >> (~&wire355)) ?
                      $signed({reg367, reg389}) : $unsigned((reg364 ?
                          reg389 : reg386))) ?
                  $unsigned($unsigned($signed(wire355))) : ((wire355[(1'h0):(1'h0)] ?
                      $unsigned(reg398) : (^reg396)) * {reg370})));
              reg402 <= $unsigned(reg370[(4'h8):(3'h7)]);
              reg403 <= reg364;
              reg404 = (reg398[(4'hf):(3'h4)] + $signed(wire356));
            end
          reg405 = {$unsigned($signed($signed((wire358 ? reg400 : reg390))))};
          for (forvar406 = (1'h0); (forvar406 < (2'h2)); forvar406 = (forvar406 + (1'h1)))
            begin
              reg407 <= $signed($unsigned($unsigned(((reg387 ?
                      reg400 : (8'hbc)) ?
                  reg396 : {wire355}))));
              reg408 <= ((({(~reg403), $unsigned(reg369)} ?
                  $unsigned((reg387 && reg389)) : $signed((reg386 ?
                      forvar406 : reg402))) ^~ $signed({(~|reg407),
                  ((8'hb8) > (8'ha3))})) - reg389[(1'h1):(1'h0)]);
              reg409 = wire356;
            end
        end
      else
        begin
          if (reg361)
            begin
              reg397 = $signed((~&$unsigned(reg398)));
            end
          else
            begin
              reg397 = $unsigned((7'h45));
            end
          reg398 <= ((forvar399[(4'he):(2'h3)] <= $signed($unsigned($unsigned(wire355)))) ?
              {$unsigned($signed((8'ha1))),
                  $unsigned($signed((wire357 ?
                      wire358 : reg400)))} : $unsigned((+(7'h48))));
          for (forvar399 = (1'h0); (forvar399 < (1'h0)); forvar399 = (forvar399 + (1'h1)))
            begin
              reg400 = reg386;
              reg401 <= {reg384};
              reg404 = $signed($signed((({reg389} ?
                  $unsigned((7'h48)) : ((8'ha0) ?
                      reg408 : reg381)) > {$unsigned(reg400), reg409})));
            end
          for (forvar405 = (1'h0); (forvar405 < (1'h1)); forvar405 = (forvar405 + (1'h1)))
            begin
              reg406 = wire355;
              reg407 <= reg369;
              reg409 = (((|(^~(~&reg402))) ?
                  (8'hbc) : (reg407[(2'h3):(1'h1)] - reg404)) || $unsigned((7'h49)));
            end
        end
      for (forvar410 = (1'h0); (forvar410 < (1'h1)); forvar410 = (forvar410 + (1'h1)))
        begin
          for (forvar411 = (1'h0); (forvar411 < (1'h0)); forvar411 = (forvar411 + (1'h1)))
            begin
              reg412 <= reg369;
            end
          for (forvar413 = (1'h0); (forvar413 < (2'h3)); forvar413 = (forvar413 + (1'h1)))
            begin
              reg414 = ((~|($unsigned({forvar397}) ?
                  forvar397[(5'h11):(3'h5)] : (&$unsigned((7'h49))))) ~^ reg409[(2'h3):(2'h2)]);
              reg415 = $signed(($signed((8'ha0)) & reg397[(3'h4):(3'h4)]));
              reg416 <= $signed((+((reg407[(1'h0):(1'h0)] >> forvar399[(5'h11):(4'hd)]) >>> $unsigned($unsigned(reg405)))));
              reg417 <= (reg415[(3'h7):(3'h4)] >> $unsigned(wire354));
              reg418 <= (reg398[(4'h8):(1'h1)] | ((wire355[(2'h2):(2'h2)] - ((~&reg402) + reg415[(2'h3):(2'h2)])) <= $unsigned((^reg387))));
            end
          for (forvar419 = (1'h0); (forvar419 < (2'h2)); forvar419 = (forvar419 + (1'h1)))
            begin
              reg420 = ((&(^(!(~|reg379)))) || (~|forvar410));
              reg421 <= wire356[(4'h9):(1'h1)];
            end
          for (forvar422 = (1'h0); (forvar422 < (2'h3)); forvar422 = (forvar422 + (1'h1)))
            begin
              reg423 <= (forvar411[(3'h4):(3'h4)] & $unsigned(($signed({forvar422,
                      forvar413}) ?
                  ($unsigned(reg390) ?
                      (reg379 >> forvar397) : reg400[(1'h0):(1'h0)]) : (^~reg384[(1'h1):(1'h0)]))));
              reg424 <= $signed(reg398[(5'h10):(4'ha)]);
            end
          for (forvar425 = (1'h0); (forvar425 < (2'h3)); forvar425 = (forvar425 + (1'h1)))
            begin
              reg426 <= $signed($signed(reg416[(3'h6):(2'h2)]));
              reg427 = reg370;
              reg428 <= ($signed(reg420) & (+{(&reg403)}));
            end
        end
    end
  always
    @(posedge clk) begin
      reg429 = reg369[(2'h3):(1'h0)];
      reg430 <= {(^~wire357[(1'h0):(1'h0)]),
          (reg381[(4'hc):(3'h5)] ?
              ((((8'haa) | reg364) ? (^~reg387) : (~&wire356)) * (^~(reg421 ?
                  wire358 : reg390))) : {reg360, $signed($signed(reg417))})};
    end
  always
    @(posedge clk) begin
      if ($signed({reg367}))
        begin
          reg431 <= (~|wire356[(3'h5):(3'h5)]);
          reg432 = {reg360[(2'h2):(2'h2)]};
          reg433 <= reg401;
          reg434 = ({((reg390[(1'h0):(1'h0)] ?
                          reg386[(4'h8):(2'h2)] : {reg421}) ?
                      $signed({reg361, wire354}) : reg364[(4'hc):(1'h0)]),
                  $unsigned($unsigned($signed(reg401)))} ?
              (8'ha0) : $signed((^~$unsigned((reg370 != (8'hb7))))));
          if (reg428[(3'h5):(1'h1)])
            begin
              reg435 <= (!reg401[(3'h4):(1'h1)]);
              reg436 = ({{reg403[(2'h2):(2'h2)], (-(-reg426))}} ?
                  $signed(reg361[(4'h8):(3'h4)]) : reg381[(4'hc):(3'h4)]);
            end
          else
            begin
              reg436 = $signed(reg417[(5'h13):(4'he)]);
              reg437 = (8'h9e);
              reg438 = $unsigned(($unsigned(wire356[(3'h7):(2'h3)]) || reg421[(4'hc):(4'hb)]));
            end
        end
      else
        begin
          reg431 <= ($signed((reg379[(4'hd):(4'h8)] & ((reg402 ~^ reg390) ?
                  $signed(reg364) : {reg367}))) ?
              reg360 : ($signed(reg434[(4'ha):(1'h0)]) + $unsigned((reg421[(2'h2):(1'h0)] == (reg434 > (8'hb1))))));
          reg433 <= (reg436 >>> reg401[(4'h8):(3'h4)]);
        end
      if (reg381)
        begin
          reg439 = $unsigned((8'hb6));
          reg440 <= $unsigned((reg430[(2'h2):(1'h0)] ^~ (((reg386 <<< reg436) > {(8'hb2),
              reg364}) >>> $signed((^~wire355)))));
          reg441 = reg396[(3'h6):(2'h2)];
          reg442 <= ((wire357[(2'h2):(2'h2)] > reg360[(2'h3):(1'h0)]) && (^~(reg412 ?
              wire358[(2'h2):(1'h0)] : ($signed(reg438) == (reg434 ?
                  wire357 : (8'h9f))))));
          reg443 <= $signed(reg403[(2'h2):(2'h2)]);
        end
      else
        begin
          if ((+reg423[(2'h2):(1'h0)]))
            begin
              reg440 <= $signed(reg423);
              reg441 = (~&$unsigned(reg402[(4'h9):(4'h9)]));
              reg442 <= reg417;
              reg443 <= (($unsigned(wire356[(4'hf):(3'h6)]) & reg396[(2'h2):(1'h0)]) >>> (reg390 >= (^~$unsigned(reg381))));
              reg444 = (!reg437);
            end
          else
            begin
              reg440 <= ({(7'h49)} ?
                  $signed($unsigned($signed(((8'hac) ?
                      (8'hac) : reg428)))) : {wire357[(1'h0):(1'h0)],
                      ($signed(reg431) <<< ((reg381 ? reg396 : reg387) ?
                          $unsigned(reg398) : $unsigned(wire356)))});
              reg441 = reg395[(2'h2):(2'h2)];
              reg442 <= $signed(reg424);
            end
          reg445 = reg367[(2'h2):(2'h2)];
          reg446 <= $unsigned((reg440 ?
              {$signed({(8'h9d), reg433}),
                  reg435} : ($unsigned({reg443}) || (|reg416))));
          if ({reg367[(2'h3):(1'h1)],
              $unsigned($signed(($signed(reg390) ?
                  $unsigned((8'hab)) : {reg434})))})
            begin
              reg447 = reg443[(2'h2):(1'h1)];
              reg448 = reg395[(2'h2):(1'h1)];
              reg449 <= reg445[(2'h2):(1'h1)];
            end
          else
            begin
              reg447 = reg444[(4'ha):(2'h3)];
              reg449 <= ({reg364[(3'h5):(1'h0)],
                  $signed(wire357[(1'h0):(1'h0)])} || $signed($unsigned($signed((reg412 ?
                  reg433 : reg444)))));
              reg450 = ($unsigned({(-((8'hb3) ? reg428 : reg445))}) ?
                  reg395 : ((wire358 ? $signed((reg444 < reg360)) : reg379) ?
                      ((|$signed(reg407)) ?
                          reg428[(2'h3):(1'h0)] : $signed(reg444[(4'h9):(1'h1)])) : (reg436 ^ (&$signed(reg426)))));
            end
        end
    end
  assign wire451 = (reg421 - reg435);
  assign wire452 = {$unsigned($signed($signed({reg412, reg440}))),
                       (~&$signed((+{(8'h9d), reg398})))};
  always
    @(posedge clk) begin
      for (forvar453 = (1'h0); (forvar453 < (1'h1)); forvar453 = (forvar453 + (1'h1)))
        begin
          reg454 = ((reg421[(5'h14):(4'ha)] ?
                  reg381[(1'h1):(1'h1)] : {$unsigned((!wire355)), {reg440}}) ?
              reg412[(4'hd):(3'h4)] : reg418);
          for (forvar455 = (1'h0); (forvar455 < (2'h3)); forvar455 = (forvar455 + (1'h1)))
            begin
              reg456 = wire354;
              reg457 <= (~^reg426);
            end
          for (forvar458 = (1'h0); (forvar458 < (1'h0)); forvar458 = (forvar458 + (1'h1)))
            begin
              reg459 = (~|reg442);
              reg460 <= $unsigned(((8'hbe) ?
                  {reg456, $unsigned((~&reg426))} : (&(~^((7'h46) < reg426)))));
            end
          reg461 = {reg360};
          reg462 <= ($signed((!$signed((reg418 ? reg435 : (7'h40))))) ?
              $unsigned(((((8'haf) ? reg398 : wire377) + (8'hbb)) ?
                  (&(reg387 ^~ (8'ha4))) : reg407[(2'h2):(1'h0)])) : $unsigned($unsigned($signed($signed(reg390)))));
        end
      reg463 = (~$signed((^$unsigned($signed(reg462)))));
      reg464 <= ({reg462,
              ((8'hab) ?
                  (forvar453 && (reg403 ?
                      (8'hb0) : reg361)) : ($signed(reg457) ?
                      $unsigned(reg379) : {forvar458, wire356}))} ?
          {wire377,
              ((reg403 <= $unsigned((8'had))) && $signed($signed((8'hb0))))} : $unsigned($signed((reg418 ?
              (reg461 ? reg433 : reg460) : reg416[(4'h8):(3'h4)]))));
      reg465 <= reg464[(3'h7):(2'h2)];
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module36
#(parameter param307 = {{(8'hbd), {{((8'hab) || (8'haa))}}}})
(y, clk, wire41, wire40, wire39, wire38, wire37);
  output wire [(32'hdd0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire41;
  input wire [(3'h4):(1'h0)] wire40;
  input wire [(5'h16):(1'h0)] wire39;
  input wire signed [(4'ha):(1'h0)] wire38;
  input wire signed [(4'hf):(1'h0)] wire37;
  wire [(4'ha):(1'h0)] wire291;
  wire signed [(4'hc):(1'h0)] wire242;
  wire signed [(3'h7):(1'h0)] wire158;
  wire [(4'hb):(1'h0)] wire140;
  wire [(4'hf):(1'h0)] wire135;
  wire signed [(4'hf):(1'h0)] wire42;
  reg signed [(3'h5):(1'h0)] reg306 = (1'h0);
  reg [(3'h5):(1'h0)] reg298 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg305 = (1'h0);
  reg [(2'h2):(1'h0)] reg302 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg301 = (1'h0);
  reg signed [(4'he):(1'h0)] reg294 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg293 = (1'h0);
  reg [(5'h11):(1'h0)] reg292 = (1'h0);
  reg [(3'h6):(1'h0)] reg285 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg282 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg278 = (1'h0);
  reg [(4'hb):(1'h0)] reg277 = (1'h0);
  reg [(5'h18):(1'h0)] reg276 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg275 = (1'h0);
  reg [(3'h5):(1'h0)] reg273 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg272 = (1'h0);
  reg [(4'h9):(1'h0)] reg271 = (1'h0);
  reg [(4'ha):(1'h0)] reg268 = (1'h0);
  reg [(2'h3):(1'h0)] reg267 = (1'h0);
  reg [(5'h16):(1'h0)] reg265 = (1'h0);
  reg [(4'hb):(1'h0)] reg264 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg261 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg260 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg258 = (1'h0);
  reg [(5'h12):(1'h0)] reg257 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg246 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg244 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg243 = (1'h0);
  reg [(5'h16):(1'h0)] reg241 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg240 = (1'h0);
  reg [(4'hd):(1'h0)] reg236 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg234 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg233 = (1'h0);
  reg [(4'ha):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg229 = (1'h0);
  reg [(5'h10):(1'h0)] reg228 = (1'h0);
  reg [(4'hf):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg224 = (1'h0);
  reg [(5'h12):(1'h0)] reg223 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg222 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg219 = (1'h0);
  reg [(3'h6):(1'h0)] reg218 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg216 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg215 = (1'h0);
  reg [(5'h14):(1'h0)] reg214 = (1'h0);
  reg [(5'h13):(1'h0)] reg211 = (1'h0);
  reg [(3'h6):(1'h0)] reg209 = (1'h0);
  reg [(4'h9):(1'h0)] reg208 = (1'h0);
  reg [(4'hd):(1'h0)] reg205 = (1'h0);
  reg [(4'hb):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg202 = (1'h0);
  reg [(5'h10):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg196 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg190 = (1'h0);
  reg signed [(4'he):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg185 = (1'h0);
  reg [(4'h9):(1'h0)] reg183 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg178 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg175 = (1'h0);
  reg [(2'h3):(1'h0)] reg172 = (1'h0);
  reg [(4'h9):(1'h0)] reg171 = (1'h0);
  reg [(5'h16):(1'h0)] reg169 = (1'h0);
  reg [(3'h5):(1'h0)] reg167 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg166 = (1'h0);
  reg [(5'h17):(1'h0)] reg165 = (1'h0);
  reg [(3'h5):(1'h0)] reg156 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg154 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg146 = (1'h0);
  reg [(5'h10):(1'h0)] reg145 = (1'h0);
  reg [(5'h10):(1'h0)] reg142 = (1'h0);
  reg [(2'h2):(1'h0)] reg139 = (1'h0);
  reg [(4'ha):(1'h0)] reg136 = (1'h0);
  reg [(5'h10):(1'h0)] reg133 = (1'h0);
  reg [(5'h14):(1'h0)] reg131 = (1'h0);
  reg [(2'h2):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg123 = (1'h0);
  reg [(2'h2):(1'h0)] reg120 = (1'h0);
  reg [(5'h18):(1'h0)] reg118 = (1'h0);
  reg [(5'h16):(1'h0)] reg117 = (1'h0);
  reg [(4'hf):(1'h0)] reg110 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg109 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg107 = (1'h0);
  reg [(5'h10):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg100 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg99 = (1'h0);
  reg [(5'h14):(1'h0)] reg98 = (1'h0);
  reg [(2'h2):(1'h0)] reg96 = (1'h0);
  reg [(2'h2):(1'h0)] reg93 = (1'h0);
  reg [(4'h8):(1'h0)] reg90 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg85 = (1'h0);
  reg [(3'h6):(1'h0)] reg84 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg79 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg77 = (1'h0);
  reg [(2'h2):(1'h0)] reg75 = (1'h0);
  reg [(4'ha):(1'h0)] reg74 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg72 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg69 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg68 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg64 = (1'h0);
  reg [(5'h10):(1'h0)] reg56 = (1'h0);
  reg [(4'h8):(1'h0)] reg55 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg52 = (1'h0);
  reg [(5'h17):(1'h0)] reg51 = (1'h0);
  reg [(4'hc):(1'h0)] reg49 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg46 = (1'h0);
  reg [(4'h9):(1'h0)] forvar304 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg300 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg299 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar298 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg297 = (1'h0);
  reg [(4'ha):(1'h0)] reg296 = (1'h0);
  reg [(5'h18):(1'h0)] reg295 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg290 = (1'h0);
  reg [(5'h12):(1'h0)] reg289 = (1'h0);
  reg [(5'h17):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar287 = (1'h0);
  reg [(4'hc):(1'h0)] reg286 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg284 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg283 = (1'h0);
  reg [(4'hc):(1'h0)] reg281 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg280 = (1'h0);
  reg [(4'hc):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg274 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar271 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg270 = (1'h0);
  reg [(3'h7):(1'h0)] reg269 = (1'h0);
  reg [(5'h16):(1'h0)] forvar266 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg263 = (1'h0);
  reg [(3'h5):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg259 = (1'h0);
  reg [(3'h6):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar254 = (1'h0);
  reg [(4'h9):(1'h0)] reg253 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg252 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg251 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg248 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar247 = (1'h0);
  reg [(3'h6):(1'h0)] forvar245 = (1'h0);
  reg [(4'hc):(1'h0)] reg239 = (1'h0);
  reg [(5'h11):(1'h0)] reg238 = (1'h0);
  reg [(4'hd):(1'h0)] reg237 = (1'h0);
  reg [(4'he):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg232 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg231 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg225 = (1'h0);
  reg signed [(4'he):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg221 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar220 = (1'h0);
  reg [(4'ha):(1'h0)] reg217 = (1'h0);
  reg [(5'h16):(1'h0)] reg213 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg212 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar207 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg206 = (1'h0);
  reg [(2'h3):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar201 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar200 = (1'h0);
  reg [(5'h12):(1'h0)] reg199 = (1'h0);
  reg [(5'h11):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg182 = (1'h0);
  reg [(5'h17):(1'h0)] reg197 = (1'h0);
  reg [(4'hd):(1'h0)] reg195 = (1'h0);
  reg [(4'hf):(1'h0)] reg194 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar193 = (1'h0);
  reg [(3'h5):(1'h0)] reg191 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg189 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg188 = (1'h0);
  reg [(2'h3):(1'h0)] reg187 = (1'h0);
  reg [(4'hb):(1'h0)] forvar184 = (1'h0);
  reg [(3'h4):(1'h0)] forvar182 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg181 = (1'h0);
  reg [(3'h4):(1'h0)] reg180 = (1'h0);
  reg [(2'h2):(1'h0)] reg179 = (1'h0);
  reg [(5'h18):(1'h0)] reg177 = (1'h0);
  reg [(2'h3):(1'h0)] reg176 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg174 = (1'h0);
  reg [(5'h17):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg170 = (1'h0);
  reg [(2'h2):(1'h0)] reg168 = (1'h0);
  reg signed [(4'he):(1'h0)] reg164 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar163 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg162 = (1'h0);
  reg [(5'h17):(1'h0)] reg161 = (1'h0);
  reg [(2'h2):(1'h0)] reg160 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg159 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar155 = (1'h0);
  reg [(4'hd):(1'h0)] reg152 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar151 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg150 = (1'h0);
  reg [(4'hd):(1'h0)] forvar149 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg148 = (1'h0);
  reg [(4'ha):(1'h0)] reg147 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg143 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar141 = (1'h0);
  reg [(4'ha):(1'h0)] reg138 = (1'h0);
  reg [(4'he):(1'h0)] forvar137 = (1'h0);
  reg [(5'h13):(1'h0)] reg134 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg132 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg130 = (1'h0);
  reg [(4'hf):(1'h0)] reg129 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg127 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg125 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg124 = (1'h0);
  reg [(4'ha):(1'h0)] forvar122 = (1'h0);
  reg [(5'h13):(1'h0)] reg121 = (1'h0);
  reg [(5'h10):(1'h0)] forvar119 = (1'h0);
  reg [(5'h17):(1'h0)] reg116 = (1'h0);
  reg [(3'h4):(1'h0)] reg115 = (1'h0);
  reg [(4'hc):(1'h0)] reg114 = (1'h0);
  reg [(5'h12):(1'h0)] forvar113 = (1'h0);
  reg [(3'h7):(1'h0)] forvar112 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg111 = (1'h0);
  reg [(4'h9):(1'h0)] reg108 = (1'h0);
  reg [(4'hc):(1'h0)] forvar106 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg105 = (1'h0);
  reg [(2'h3):(1'h0)] forvar103 = (1'h0);
  reg [(5'h12):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg101 = (1'h0);
  reg [(4'hc):(1'h0)] forvar97 = (1'h0);
  reg [(4'hf):(1'h0)] reg95 = (1'h0);
  reg [(3'h7):(1'h0)] reg94 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg92 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg91 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg88 = (1'h0);
  reg [(2'h2):(1'h0)] reg87 = (1'h0);
  reg [(4'h9):(1'h0)] reg86 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg83 = (1'h0);
  reg [(2'h2):(1'h0)] reg82 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg81 = (1'h0);
  reg [(3'h6):(1'h0)] forvar78 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg73 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar72 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg71 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg70 = (1'h0);
  reg [(5'h18):(1'h0)] forvar67 = (1'h0);
  reg [(5'h18):(1'h0)] reg66 = (1'h0);
  reg [(5'h10):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg63 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg62 = (1'h0);
  reg [(5'h12):(1'h0)] reg61 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg60 = (1'h0);
  reg [(5'h13):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar58 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg57 = (1'h0);
  reg [(4'hd):(1'h0)] reg54 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg53 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar50 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg48 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg47 = (1'h0);
  reg [(5'h11):(1'h0)] forvar44 = (1'h0);
  reg [(3'h6):(1'h0)] reg43 = (1'h0);
  reg [(4'ha):(1'h0)] reg45 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg44 = (1'h0);
  reg [(5'h13):(1'h0)] forvar43 = (1'h0);
  assign y = {wire291,
                 wire242,
                 wire158,
                 wire140,
                 wire135,
                 wire42,
                 reg306,
                 reg298,
                 reg305,
                 reg302,
                 reg301,
                 reg294,
                 reg293,
                 reg292,
                 reg285,
                 reg282,
                 reg278,
                 reg277,
                 reg276,
                 reg275,
                 reg273,
                 reg272,
                 reg271,
                 reg268,
                 reg267,
                 reg265,
                 reg264,
                 reg261,
                 reg260,
                 reg258,
                 reg257,
                 reg255,
                 reg250,
                 reg246,
                 reg244,
                 reg243,
                 reg241,
                 reg240,
                 reg236,
                 reg234,
                 reg233,
                 reg230,
                 reg229,
                 reg228,
                 reg226,
                 reg224,
                 reg223,
                 reg222,
                 reg219,
                 reg218,
                 reg216,
                 reg215,
                 reg214,
                 reg211,
                 reg209,
                 reg208,
                 reg205,
                 reg203,
                 reg202,
                 reg198,
                 reg196,
                 reg192,
                 reg190,
                 reg186,
                 reg185,
                 reg183,
                 reg178,
                 reg175,
                 reg172,
                 reg171,
                 reg169,
                 reg167,
                 reg166,
                 reg165,
                 reg156,
                 reg154,
                 reg153,
                 reg146,
                 reg145,
                 reg142,
                 reg139,
                 reg136,
                 reg133,
                 reg131,
                 reg128,
                 reg126,
                 reg123,
                 reg120,
                 reg118,
                 reg117,
                 reg110,
                 reg109,
                 reg107,
                 reg104,
                 reg100,
                 reg99,
                 reg98,
                 reg96,
                 reg93,
                 reg90,
                 reg89,
                 reg85,
                 reg84,
                 reg80,
                 reg79,
                 reg77,
                 reg75,
                 reg74,
                 reg72,
                 reg69,
                 reg68,
                 reg64,
                 reg56,
                 reg55,
                 reg52,
                 reg51,
                 reg49,
                 reg46,
                 forvar304,
                 reg303,
                 reg300,
                 reg299,
                 forvar298,
                 reg297,
                 reg296,
                 reg295,
                 reg290,
                 reg289,
                 reg288,
                 forvar287,
                 reg286,
                 reg284,
                 reg283,
                 reg281,
                 reg280,
                 reg279,
                 reg274,
                 forvar271,
                 reg270,
                 reg269,
                 forvar266,
                 reg263,
                 reg262,
                 reg259,
                 reg256,
                 forvar254,
                 reg253,
                 reg252,
                 reg251,
                 reg249,
                 reg248,
                 forvar247,
                 forvar245,
                 reg239,
                 reg238,
                 reg237,
                 reg235,
                 reg232,
                 reg231,
                 reg227,
                 reg225,
                 reg220,
                 reg221,
                 forvar220,
                 reg217,
                 reg213,
                 reg212,
                 reg210,
                 forvar207,
                 reg206,
                 reg204,
                 forvar201,
                 forvar200,
                 reg199,
                 reg184,
                 reg182,
                 reg197,
                 reg195,
                 reg194,
                 forvar193,
                 reg191,
                 reg189,
                 reg188,
                 reg187,
                 forvar184,
                 forvar182,
                 reg181,
                 reg180,
                 reg179,
                 reg177,
                 reg176,
                 reg174,
                 reg173,
                 reg170,
                 reg168,
                 reg164,
                 forvar163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg157,
                 forvar155,
                 reg152,
                 forvar151,
                 reg150,
                 forvar149,
                 reg148,
                 reg147,
                 reg144,
                 reg143,
                 forvar141,
                 reg138,
                 forvar137,
                 reg134,
                 reg132,
                 reg130,
                 reg129,
                 reg127,
                 reg125,
                 reg124,
                 forvar122,
                 reg121,
                 forvar119,
                 reg116,
                 reg115,
                 reg114,
                 forvar113,
                 forvar112,
                 reg111,
                 reg108,
                 forvar106,
                 reg105,
                 forvar103,
                 reg102,
                 reg101,
                 forvar97,
                 reg95,
                 reg94,
                 reg92,
                 reg91,
                 reg88,
                 reg87,
                 reg86,
                 reg83,
                 reg82,
                 reg81,
                 forvar78,
                 reg76,
                 reg73,
                 forvar72,
                 reg71,
                 reg70,
                 forvar67,
                 reg66,
                 reg65,
                 reg63,
                 reg62,
                 reg61,
                 reg60,
                 reg59,
                 forvar58,
                 reg57,
                 reg54,
                 reg53,
                 forvar50,
                 reg48,
                 reg47,
                 forvar44,
                 reg43,
                 reg45,
                 reg44,
                 forvar43,
                 (1'h0)};
  assign wire42 = $signed($unsigned(({$signed(wire38),
                      (wire38 | wire37)} != $unsigned($unsigned((8'hbd))))));
  always
    @(posedge clk) begin
      if (wire37)
        begin
          for (forvar43 = (1'h0); (forvar43 < (1'h1)); forvar43 = (forvar43 + (1'h1)))
            begin
              reg44 = (~&(wire41 ?
                  $unsigned($unsigned((wire39 ?
                      wire39 : wire39))) : (~^wire38)));
              reg45 = wire38[(3'h4):(3'h4)];
            end
          reg46 <= wire37;
        end
      else
        begin
          reg43 = wire39[(4'ha):(4'h8)];
          for (forvar44 = (1'h0); (forvar44 < (2'h2)); forvar44 = (forvar44 + (1'h1)))
            begin
              reg45 = $unsigned(($unsigned((wire40[(3'h4):(2'h3)] ^~ wire40)) > $signed($unsigned({(7'h43)}))));
              reg47 = ($unsigned($signed(reg46)) != ((((+wire41) ?
                          (wire40 == wire40) : $unsigned(reg43)) ?
                      (&{forvar43}) : {forvar43[(4'h8):(2'h3)]}) ?
                  wire40 : ((^~(wire42 ?
                      forvar44 : forvar44)) <<< $signed({wire40, wire39}))));
              reg48 = ($unsigned($signed($signed($unsigned((8'ha2))))) ?
                  forvar44[(3'h6):(1'h0)] : reg45[(3'h4):(2'h3)]);
              reg49 <= wire38[(4'ha):(4'h8)];
            end
          for (forvar50 = (1'h0); (forvar50 < (3'h4)); forvar50 = (forvar50 + (1'h1)))
            begin
              reg51 <= reg45;
              reg52 <= ($signed(($signed(forvar50[(3'h6):(1'h0)]) + (((8'hba) < reg44) ?
                      wire38[(1'h1):(1'h1)] : wire38[(3'h7):(3'h6)]))) ?
                  $unsigned((&$signed((reg47 ?
                      wire37 : wire42)))) : (reg47 <= (reg46 ?
                      ((reg47 ^~ forvar50) ?
                          reg45[(4'h9):(4'h8)] : (forvar43 ?
                              (7'h44) : reg45)) : reg46[(1'h1):(1'h0)])));
              reg53 = (wire38 ?
                  ($signed((+$signed(wire37))) ?
                      (^{(reg43 ?
                              (7'h42) : forvar50)}) : {reg45[(2'h2):(2'h2)]}) : $signed((8'ha0)));
              reg54 = (reg52 ?
                  ($signed(((wire41 ? wire40 : (8'ha4)) ?
                          wire37[(1'h0):(1'h0)] : {wire37})) ?
                      $signed((+(wire37 ?
                          wire38 : wire40))) : (forvar43[(5'h12):(5'h11)] >> $signed((wire38 >> (8'h9f))))) : reg53[(5'h12):(4'h9)]);
              reg55 <= $signed(wire42[(3'h7):(1'h1)]);
            end
          reg56 <= {$unsigned((reg47[(3'h4):(1'h0)] || $signed((reg44 ?
                  wire42 : wire39)))),
              (~(!forvar43[(4'he):(3'h4)]))};
          reg57 = (forvar44[(2'h2):(1'h0)] >= $unsigned({$signed($signed(forvar50))}));
        end
      for (forvar58 = (1'h0); (forvar58 < (2'h2)); forvar58 = (forvar58 + (1'h1)))
        begin
          if ((-wire42))
            begin
              reg59 = $signed(forvar58[(4'ha):(2'h3)]);
              reg60 = {(8'ha9), $signed(forvar58)};
              reg61 = {reg48};
              reg62 = ((($signed(reg57) ?
                      $signed($unsigned(wire41)) : reg49[(3'h4):(1'h0)]) ?
                  ({(forvar44 ? forvar44 : reg59), (|forvar50)} ?
                      (+reg59) : reg52) : $signed((~|(~^wire37)))) ~^ $unsigned((~|($signed(forvar44) & (~^reg47)))));
              reg63 = (~^$unsigned({(+$unsigned(reg47))}));
            end
          else
            begin
              reg59 = reg49;
              reg60 = (forvar43 ?
                  {(forvar50[(4'hb):(4'hb)] ^~ (^~(^~wire40)))} : $unsigned(forvar43[(4'he):(4'hb)]));
              reg64 <= (!reg54);
              reg65 = (!((~{(~&reg44), (forvar44 ~^ reg57)}) ?
                  (reg47[(1'h1):(1'h1)] <<< $unsigned(reg45)) : $signed($unsigned($signed(reg52)))));
              reg66 = (^($unsigned(((~^reg45) & ((8'hab) ?
                  reg56 : reg65))) || $unsigned((8'hb3))));
            end
          for (forvar67 = (1'h0); (forvar67 < (1'h0)); forvar67 = (forvar67 + (1'h1)))
            begin
              reg68 <= $signed(reg63[(4'he):(3'h4)]);
              reg69 <= $signed((wire40[(2'h2):(1'h1)] + $unsigned((reg62 ?
                  reg46 : $unsigned(wire42)))));
              reg70 = reg43[(3'h5):(1'h0)];
              reg71 = forvar67;
            end
        end
      if ({($unsigned($signed(reg51)) ~^ forvar67),
          {$signed(($signed(reg65) * reg49[(4'ha):(3'h7)])),
              (~(!wire41[(3'h4):(1'h1)]))}})
        begin
          reg72 <= reg71;
        end
      else
        begin
          for (forvar72 = (1'h0); (forvar72 < (3'h4)); forvar72 = (forvar72 + (1'h1)))
            begin
              reg73 = $unsigned(({reg56[(3'h6):(1'h1)], (~^reg52)} ?
                  reg72[(4'h8):(3'h5)] : (reg63 ?
                      $signed({reg64, reg43}) : {reg72})));
              reg74 <= $unsigned({(8'hb5)});
              reg75 <= wire42[(2'h2):(2'h2)];
              reg76 = (7'h40);
              reg77 <= (reg69 - (-(($signed(reg66) >= ((8'hab) ?
                      (8'hae) : reg69)) ?
                  reg60 : reg60)));
            end
          for (forvar78 = (1'h0); (forvar78 < (1'h0)); forvar78 = (forvar78 + (1'h1)))
            begin
              reg79 <= reg47;
              reg80 <= ((reg47 >> (~^($unsigned(reg57) ^~ {reg54}))) ?
                  ((reg62 ^ reg63) ?
                      (+$unsigned((forvar78 && wire40))) : (wire39[(4'hc):(3'h6)] ^~ $unsigned(reg52[(4'hd):(1'h0)]))) : (~|($signed((|reg47)) ?
                      $unsigned((reg79 ? reg71 : reg49)) : (8'ha9))));
              reg81 = wire37;
              reg82 = ($unsigned((+reg57[(4'hd):(4'ha)])) ?
                  (~&wire40) : $unsigned(reg73));
              reg83 = $signed($unsigned((reg60[(4'h9):(3'h5)] ?
                  $unsigned($unsigned(reg77)) : ((reg44 && reg51) | $unsigned(forvar58)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg84 <= {reg68[(4'h9):(2'h2)],
          ((reg77[(3'h5):(1'h1)] ?
                  (reg46 ?
                      (reg80 ? reg46 : reg56) : (reg64 ?
                          reg52 : (8'hb7))) : wire40) ?
              $signed(reg55[(2'h3):(1'h1)]) : reg74)};
    end
  always
    @(posedge clk) begin
      reg85 <= reg55;
      if ($unsigned(wire40))
        begin
          reg86 = reg69;
          reg87 = $unsigned({$signed($signed(wire38[(3'h6):(1'h1)]))});
          reg88 = ($unsigned($unsigned(reg77[(2'h2):(1'h1)])) ?
              reg79 : $unsigned(({(^reg75), (reg49 ? reg74 : (8'hbc))} ?
                  ((reg87 ? reg52 : reg87) * ((8'hbb) ?
                      (8'h9e) : reg75)) : (^~reg69[(4'hc):(2'h2)]))));
          reg89 <= $unsigned(reg75[(1'h1):(1'h1)]);
        end
      else
        begin
          if ($unsigned(reg75))
            begin
              reg89 <= $signed(reg80);
              reg90 <= (wire41 ?
                  (reg87[(2'h2):(1'h0)] * reg84[(3'h5):(1'h1)]) : {(&((reg85 <<< reg56) ?
                          (+wire39) : (!(7'h40)))),
                      reg74[(4'h8):(4'h8)]});
              reg91 = {$signed($signed(reg88[(4'hd):(4'h8)])),
                  {{((wire41 ? (7'h43) : (7'h47)) ? $signed(reg79) : wire38),
                          ((8'hba) & $unsigned(reg79))}}};
              reg92 = ((~^$unsigned(((!reg84) ?
                  $unsigned((8'ha2)) : wire39[(4'hf):(4'ha)]))) != reg72);
              reg93 <= {reg68};
            end
          else
            begin
              reg89 <= ($signed(reg86[(4'h8):(4'h8)]) < $signed($unsigned((~(&wire38)))));
              reg90 <= reg93[(2'h2):(1'h0)];
              reg91 = reg69;
            end
        end
      reg94 = wire40[(1'h0):(1'h0)];
      reg95 = (reg55 ?
          wire39[(4'h9):(4'h8)] : ((7'h43) ?
              $signed($signed({reg90})) : reg49));
    end
  always
    @(posedge clk) begin
      reg96 <= reg56;
      if (({(({wire40, reg69} ? reg64 : (reg69 - reg89)) ?
                  $signed({reg74, reg55}) : (~|(reg52 - wire40)))} ?
          $unsigned({(+reg80[(2'h2):(1'h1)]),
              (8'ha4)}) : $signed($unsigned((~&reg85)))))
        begin
          for (forvar97 = (1'h0); (forvar97 < (1'h1)); forvar97 = (forvar97 + (1'h1)))
            begin
              reg98 <= reg96[(1'h1):(1'h1)];
              reg99 <= reg80[(3'h6):(3'h6)];
              reg100 <= reg55;
              reg101 = (&wire42[(4'ha):(3'h7)]);
              reg102 = $signed(forvar97);
            end
          for (forvar103 = (1'h0); (forvar103 < (3'h4)); forvar103 = (forvar103 + (1'h1)))
            begin
              reg104 <= (($unsigned(($unsigned(reg72) ?
                      (reg100 ?
                          (8'hb8) : wire37) : forvar97[(4'hb):(1'h1)])) <<< (&($unsigned(reg75) << (+wire38)))) ?
                  ($signed($unsigned((|reg93))) ?
                      reg74 : (~|reg79)) : ($signed($signed((reg98 == reg89))) ?
                      ((~&reg69[(4'he):(4'h9)]) ?
                          $unsigned({reg75}) : $signed(wire39)) : reg84));
              reg105 = $signed($unsigned($signed((|reg79[(4'ha):(1'h0)]))));
            end
          for (forvar106 = (1'h0); (forvar106 < (2'h2)); forvar106 = (forvar106 + (1'h1)))
            begin
              reg107 <= ({reg77,
                      ($unsigned(wire39) < (reg75 * (reg101 ?
                          forvar103 : reg93)))} ?
                  {$unsigned($unsigned((^reg102))),
                      (-$unsigned(reg77))} : ((($unsigned(reg79) ?
                      (reg101 ? reg100 : reg49) : {wire42,
                          reg101}) | (~&(forvar106 >>> reg74))) > reg85[(4'hd):(3'h7)]));
              reg108 = forvar103[(1'h1):(1'h1)];
              reg109 <= $unsigned((wire42[(4'h9):(2'h2)] ?
                  (~&(-$unsigned(reg102))) : (($unsigned(reg64) * $signed(forvar103)) | (-reg101[(4'hb):(3'h5)]))));
              reg110 <= (^reg80[(3'h4):(3'h4)]);
            end
        end
      else
        begin
          for (forvar97 = (1'h0); (forvar97 < (1'h1)); forvar97 = (forvar97 + (1'h1)))
            begin
              reg98 <= reg108[(3'h7):(3'h7)];
            end
        end
      reg111 = $signed($unsigned($unsigned(($signed(reg56) ^ reg107[(3'h6):(3'h6)]))));
    end
  always
    @(posedge clk) begin
      for (forvar112 = (1'h0); (forvar112 < (3'h4)); forvar112 = (forvar112 + (1'h1)))
        begin
          for (forvar113 = (1'h0); (forvar113 < (1'h0)); forvar113 = (forvar113 + (1'h1)))
            begin
              reg114 = (~reg75);
              reg115 = $signed(reg75);
            end
          if (reg49)
            begin
              reg116 = $unsigned((reg80[(3'h7):(3'h5)] ~^ $signed((reg74 >= {reg89,
                  reg107}))));
            end
          else
            begin
              reg117 <= reg90[(2'h2):(1'h1)];
              reg118 <= {(^$signed(reg77))};
            end
          for (forvar119 = (1'h0); (forvar119 < (2'h2)); forvar119 = (forvar119 + (1'h1)))
            begin
              reg120 <= $signed(({((reg89 ~^ reg75) ?
                          $signed(reg116) : reg52[(4'hf):(4'hc)]),
                      ({reg84, wire38} ^ (~reg115))} ?
                  $signed(reg46) : ($unsigned(((8'ha4) < reg117)) ?
                      reg100 : $signed((reg93 ? reg117 : reg51)))));
              reg121 = $signed(((($signed(reg115) > (~&reg80)) ^~ $unsigned({reg120})) | ((reg72 <= $unsigned(reg107)) | $signed(reg90[(3'h4):(2'h2)]))));
            end
          for (forvar122 = (1'h0); (forvar122 < (2'h3)); forvar122 = (forvar122 + (1'h1)))
            begin
              reg123 <= (($signed($unsigned((wire42 < reg117))) != reg110) * ($signed(reg110) > $signed((((8'hbc) <<< reg104) ?
                  ((8'hb8) ? wire37 : reg69) : reg89[(3'h6):(1'h1)]))));
              reg124 = reg115;
              reg125 = reg55;
              reg126 <= (~reg72);
              reg127 = (($signed(((^~reg96) <<< $signed(forvar122))) ^~ reg89) <<< {($signed((reg85 <<< reg107)) << ((~^reg114) || $signed(reg99)))});
            end
          reg128 <= reg69[(3'h4):(1'h0)];
        end
      reg129 = reg114;
      reg130 = (~$unsigned(reg123[(3'h6):(3'h5)]));
      reg131 <= ((+($signed((~^reg123)) + $unsigned((+reg55)))) ^~ (&(((&reg118) ?
              (^~reg64) : $signed(wire37)) ?
          (reg72 ?
              $unsigned(forvar112) : $signed(reg130)) : (reg80[(3'h7):(3'h4)] ~^ reg129[(4'hf):(4'hc)]))));
    end
  always
    @(posedge clk) begin
      reg132 = wire37[(4'ha):(2'h2)];
      reg133 <= reg80[(2'h3):(1'h0)];
      reg134 = reg51[(4'hb):(4'hb)];
    end
  assign wire135 = reg46;
  always
    @(posedge clk) begin
      reg136 <= $unsigned(reg52[(5'h11):(3'h4)]);
    end
  always
    @(posedge clk) begin
      for (forvar137 = (1'h0); (forvar137 < (1'h0)); forvar137 = (forvar137 + (1'h1)))
        begin
          if ($signed($unsigned(((reg72 >> (~&reg118)) >> ($signed(reg80) ?
              (reg136 ? reg85 : reg69) : {reg110, reg49})))))
            begin
              reg138 = $unsigned(($unsigned($signed($signed(reg80))) - $unsigned(reg98)));
            end
          else
            begin
              reg139 <= reg93;
            end
        end
    end
  assign wire140 = $unsigned(wire135);
  always
    @(posedge clk) begin
      for (forvar141 = (1'h0); (forvar141 < (1'h1)); forvar141 = (forvar141 + (1'h1)))
        begin
          if (({reg77[(3'h4):(2'h3)], reg136[(3'h4):(3'h4)]} + reg128))
            begin
              reg142 <= reg98;
            end
          else
            begin
              reg143 = ((reg139[(2'h2):(2'h2)] || ((^$signed((7'h43))) << wire38)) | $signed($unsigned(((8'hb6) && (~|reg56)))));
              reg144 = (|$signed((reg85[(4'he):(3'h5)] <= {(&reg46)})));
              reg145 <= (~&$unsigned((^($signed((7'h43)) ?
                  (wire135 ? forvar141 : reg68) : $signed(reg79)))));
            end
          reg146 <= reg77;
          reg147 = wire39[(4'hf):(3'h7)];
          reg148 = (8'hb4);
        end
      for (forvar149 = (1'h0); (forvar149 < (2'h3)); forvar149 = (forvar149 + (1'h1)))
        begin
          reg150 = wire41[(1'h1):(1'h0)];
          for (forvar151 = (1'h0); (forvar151 < (1'h1)); forvar151 = (forvar151 + (1'h1)))
            begin
              reg152 = (reg64 || reg144[(1'h0):(1'h0)]);
              reg153 <= ((^~$unsigned(reg68[(3'h5):(1'h1)])) == $signed($signed($signed((reg139 <= reg145)))));
            end
          reg154 <= (^{($unsigned(((8'hb2) <= (7'h4a))) || $signed({reg98,
                  forvar151}))});
          for (forvar155 = (1'h0); (forvar155 < (1'h1)); forvar155 = (forvar155 + (1'h1)))
            begin
              reg156 <= $unsigned($signed((~^((&(8'ha8)) * (&reg128)))));
            end
        end
      reg157 = ((reg146 && reg126) <= $signed({(^~$unsigned(reg80)),
          ($unsigned(reg126) ^~ $signed(reg146))}));
    end
  assign wire158 = (reg156[(2'h2):(1'h1)] | ($unsigned($signed(wire42)) ?
                       {(~^reg145)} : (^((+reg72) ?
                           (wire40 ? reg109 : reg89) : ((8'hbe) <= (8'hbd))))));
  always
    @(posedge clk) begin
      reg159 = {$unsigned(reg84)};
      reg160 = ((-{reg120,
          (reg104[(3'h7):(3'h5)] != (|reg139))}) < $unsigned(((reg118 <= (reg52 ?
              reg126 : reg146)) ?
          (8'ha0) : wire40[(3'h4):(1'h0)])));
      reg161 = $unsigned($unsigned(wire37));
    end
  always
    @(posedge clk) begin
      reg162 = reg64[(1'h1):(1'h0)];
      for (forvar163 = (1'h0); (forvar163 < (1'h0)); forvar163 = (forvar163 + (1'h1)))
        begin
          reg164 = $signed($unsigned(reg64[(2'h3):(2'h2)]));
          if (($unsigned(reg123) * (~^(+$signed((wire140 ~^ reg98))))))
            begin
              reg165 <= $unsigned(reg117[(5'h11):(4'he)]);
              reg166 <= ({(($unsigned(reg46) && (reg52 ? reg49 : reg131)) ?
                          $unsigned(reg93[(2'h2):(2'h2)]) : $unsigned({reg156,
                              reg154})),
                      reg133[(4'hd):(2'h3)]} ?
                  reg133 : reg72[(4'h8):(3'h5)]);
              reg167 <= reg162;
              reg168 = {(~|(reg75 ?
                      ((&reg133) > (|reg146)) : {((8'hae) ?
                              reg118 : wire40)}))};
              reg169 <= $signed($signed(((^$signed(reg77)) <= $unsigned(reg166))));
            end
          else
            begin
              reg168 = ((((reg64 ? reg153[(3'h6):(1'h1)] : (&(7'h45))) ?
                  (~&(8'hb5)) : ((reg75 ^~ wire158) < (reg110 ?
                      reg167 : (8'hac)))) || (((reg142 <= wire158) >> (reg118 ?
                  (8'ha8) : forvar163)) ^ {reg69[(4'h9):(3'h5)],
                  $unsigned(reg51)})) || (^(reg131[(5'h10):(4'hd)] ?
                  wire42[(3'h6):(3'h4)] : reg93)));
            end
          if (reg69[(4'h8):(3'h5)])
            begin
              reg170 = reg169;
              reg171 <= (^~({$signed(reg46[(3'h4):(2'h3)]),
                  reg110} && ((wire42[(1'h1):(1'h0)] + (wire39 ?
                  reg128 : wire140)) ~^ $signed({reg46, reg69}))));
              reg172 <= (8'hbf);
              reg173 = reg120;
            end
          else
            begin
              reg171 <= $unsigned(reg123);
              reg172 <= ((8'h9f) ^ ((&$signed(((8'haa) ? reg99 : (8'hac)))) ?
                  {(reg52 ? $signed(reg154) : {reg72, reg136}),
                      (reg84[(2'h3):(2'h3)] << reg164[(3'h4):(1'h0)])} : (~$unsigned($unsigned(reg156)))));
            end
          reg174 = reg84;
          if (wire39[(2'h3):(1'h0)])
            begin
              reg175 <= (8'had);
              reg176 = $unsigned($signed($signed((-reg154[(4'hc):(1'h0)]))));
              reg177 = $unsigned(wire40[(1'h1):(1'h0)]);
              reg178 <= {reg52};
            end
          else
            begin
              reg175 <= (&{{((reg165 ~^ reg84) ?
                          (reg75 ? reg146 : reg178) : $signed(wire158)),
                      ($unsigned(reg79) << (reg85 ? reg98 : reg168))}});
              reg178 <= reg84;
              reg179 = (^reg120[(1'h0):(1'h0)]);
              reg180 = ({(^(|reg170))} ?
                  ({{reg174[(3'h4):(1'h0)],
                          (reg46 <= wire40)}} >= ($unsigned((reg49 ?
                      (7'h41) : wire41)) | ((reg46 ? wire37 : reg69) ?
                      $signed((8'hb7)) : (reg120 ?
                          reg93 : reg131)))) : reg104[(2'h2):(1'h0)]);
            end
        end
      reg181 = {($unsigned($signed((~^reg168))) ?
              $unsigned({(reg107 >>> (8'hbc))}) : ((~&$signed(reg165)) ?
                  (|((8'hb0) ? reg96 : reg98)) : (~|reg84))),
          ($unsigned($unsigned($unsigned(reg85))) ?
              reg178[(4'h9):(2'h3)] : $unsigned($signed($unsigned(reg120))))};
      if (reg77)
        begin
          for (forvar182 = (1'h0); (forvar182 < (2'h3)); forvar182 = (forvar182 + (1'h1)))
            begin
              reg183 <= (~&reg153);
            end
          for (forvar184 = (1'h0); (forvar184 < (2'h3)); forvar184 = (forvar184 + (1'h1)))
            begin
              reg185 <= reg179[(1'h0):(1'h0)];
              reg186 <= reg51;
              reg187 = (reg178 <= reg89[(4'h8):(2'h3)]);
              reg188 = (reg169[(5'h10):(3'h4)] >= reg79);
              reg189 = reg131;
            end
          if ((^(($signed((reg110 >> reg179)) ?
              (reg176[(2'h3):(1'h0)] * reg171) : (+{reg164,
                  wire41})) * (reg79[(2'h2):(1'h0)] ?
              $unsigned($signed(wire39)) : $signed($signed(reg133))))))
            begin
              reg190 <= $unsigned($unsigned(reg185));
              reg191 = $signed((($unsigned((reg165 ?
                      reg153 : reg80)) & {$signed(wire140)}) ?
                  {reg49[(4'h8):(1'h1)],
                      reg126[(2'h2):(1'h0)]} : $unsigned(reg142[(4'h8):(1'h0)])));
            end
          else
            begin
              reg190 <= reg96[(1'h1):(1'h0)];
              reg191 = wire40[(3'h4):(1'h0)];
            end
          reg192 <= reg165[(3'h6):(1'h1)];
          for (forvar193 = (1'h0); (forvar193 < (1'h0)); forvar193 = (forvar193 + (1'h1)))
            begin
              reg194 = {{reg89[(2'h2):(2'h2)]}, ($signed(reg139) | reg110)};
              reg195 = reg186[(3'h5):(1'h0)];
              reg196 <= reg118;
              reg197 = $unsigned((|(((^~reg181) >= (reg177 ? reg77 : (8'hbd))) ?
                  $unsigned($signed((8'hb3))) : $signed((-reg55)))));
              reg198 <= (~reg162);
            end
        end
      else
        begin
          reg182 = $unsigned((reg180 << reg131[(4'hf):(3'h4)]));
          reg183 <= {$unsigned(wire37), (^~$signed({reg188[(3'h6):(1'h0)]}))};
          if (((!$signed($signed($signed(reg100)))) <= $signed(reg171[(2'h2):(1'h1)])))
            begin
              reg184 = $signed($unsigned((reg110 >= (+reg110[(4'hd):(4'h9)]))));
              reg187 = ((((~&reg74[(1'h1):(1'h1)]) ?
                          reg139[(1'h0):(1'h0)] : reg188[(2'h3):(1'h0)]) ?
                      $unsigned($unsigned(reg123)) : (reg164[(3'h6):(2'h2)] ?
                          (((7'h45) >= reg142) ?
                              (~|(8'hb2)) : $unsigned(reg174)) : ($unsigned(reg51) ?
                              (-reg191) : $signed(reg117)))) ?
                  reg100 : reg72[(3'h7):(3'h7)]);
              reg188 = ((~reg100[(2'h3):(2'h3)]) ?
                  reg68 : $unsigned((reg196[(4'he):(2'h2)] ?
                      {(reg128 * reg153),
                          (wire38 ? reg89 : reg197)} : ((reg128 != reg74) ?
                          $unsigned(reg46) : $signed(reg90)))));
              reg189 = reg46[(1'h1):(1'h0)];
              reg191 = (+reg98);
            end
          else
            begin
              reg185 <= $unsigned(({(reg175 ?
                          (reg128 ? reg104 : reg185) : $signed((8'ha6))),
                      forvar163[(3'h5):(1'h1)]} ?
                  (-(!(reg186 ~^ reg72))) : reg118));
            end
        end
    end
  always
    @(posedge clk) begin
      reg199 = $unsigned($unsigned({({reg74} + $unsigned(reg85))}));
      for (forvar200 = (1'h0); (forvar200 < (3'h4)); forvar200 = (forvar200 + (1'h1)))
        begin
          for (forvar201 = (1'h0); (forvar201 < (3'h4)); forvar201 = (forvar201 + (1'h1)))
            begin
              reg202 <= $signed((reg74 ? reg118 : $signed(reg185)));
              reg203 <= ($signed((~^$unsigned(reg52))) ~^ $unsigned(reg98[(4'hf):(4'hc)]));
              reg204 = (reg190 <= $unsigned(reg139[(1'h1):(1'h1)]));
              reg205 <= (reg99[(5'h17):(5'h12)] << $signed($signed((reg89 ?
                  reg199[(4'hc):(4'h9)] : reg49[(3'h5):(1'h0)]))));
            end
          reg206 = reg99;
          for (forvar207 = (1'h0); (forvar207 < (1'h0)); forvar207 = (forvar207 + (1'h1)))
            begin
              reg208 <= (($unsigned($unsigned($signed(reg109))) ^~ reg202[(5'h15):(5'h14)]) ?
                  reg117 : $unsigned($unsigned({(reg205 ? reg96 : wire40),
                      reg46[(2'h3):(2'h2)]})));
            end
          if ((~|((((reg133 ? (8'h9f) : reg79) < (reg192 ^~ reg131)) ?
                  (!(reg186 ? reg77 : reg204)) : $signed((8'h9c))) ?
              (~{{reg89, reg128}, (reg185 > reg156)}) : reg183)))
            begin
              reg209 <= (($unsigned((~|{reg90})) < (((reg90 ^ reg46) > (~&reg123)) <= reg104)) || ($signed($unsigned($signed(reg146))) ?
                  ((8'hb6) ?
                      ((&reg100) ^~ (^~wire158)) : (-reg146[(3'h5):(1'h0)])) : (reg96 - wire40)));
              reg210 = (8'haa);
              reg211 <= ((8'h9d) ? (!reg80[(4'ha):(3'h5)]) : wire135);
              reg212 = $signed((reg136[(4'h9):(4'h8)] ?
                  $unsigned(({reg104,
                      reg153} << $unsigned(wire38))) : reg203[(1'h0):(1'h0)]));
            end
          else
            begin
              reg209 <= wire39[(4'h8):(3'h5)];
            end
          reg213 = reg153;
        end
      if ((^$signed(reg96)))
        begin
          if ($unsigned($signed(((8'hbf) ?
              $unsigned(reg172[(1'h1):(1'h1)]) : $signed((reg72 ?
                  reg156 : reg192))))))
            begin
              reg214 <= (-$unsigned($unsigned(({reg46} * $signed(reg172)))));
            end
          else
            begin
              reg214 <= reg104[(1'h0):(1'h0)];
              reg215 <= reg210;
              reg216 <= $unsigned(reg96);
            end
          reg217 = reg216;
          reg218 <= ($unsigned({((reg72 & reg80) ?
                      reg55[(3'h4):(3'h4)] : (!reg209))}) ?
              reg49[(4'hb):(2'h3)] : $unsigned($signed($unsigned({forvar201,
                  reg190}))));
          reg219 <= $unsigned(reg64);
          for (forvar220 = (1'h0); (forvar220 < (2'h3)); forvar220 = (forvar220 + (1'h1)))
            begin
              reg221 = ({$unsigned((reg154 ~^ {reg46}))} ?
                  (reg136 ?
                      $unsigned($signed($signed(reg217))) : ((&(reg139 ?
                          reg109 : reg136)) ^ ((^~reg85) ~^ $unsigned(reg172)))) : ((^~$unsigned((^~reg146))) + $unsigned(((reg196 ?
                      reg75 : reg208) < (reg110 ? reg99 : reg79)))));
              reg222 <= $signed(reg100);
              reg223 <= (+reg219[(3'h7):(2'h2)]);
              reg224 <= wire37;
            end
        end
      else
        begin
          if ((reg68 * $unsigned($unsigned((!{reg107})))))
            begin
              reg217 = $unsigned(((($unsigned(reg153) ^~ ((8'hb0) >>> (8'hb8))) >> reg55[(1'h0):(1'h0)]) ?
                  (~{(|(8'ha1))}) : reg120[(1'h0):(1'h0)]));
            end
          else
            begin
              reg214 <= reg221;
              reg217 = (+reg167);
              reg220 = (reg175 ?
                  $signed(($signed(reg80[(2'h2):(2'h2)]) ?
                      ($signed(reg90) && (reg90 ?
                          reg90 : reg100)) : reg210[(4'he):(3'h4)])) : {reg154,
                      $unsigned(($signed(reg74) * (reg85 - reg64)))});
              reg222 <= {$unsigned($unsigned(reg216[(4'h8):(3'h4)])),
                  $unsigned($signed((+(reg77 & reg69))))};
              reg225 = (((reg64[(2'h3):(1'h0)] ?
                  ($signed(reg117) < (~forvar207)) : ($unsigned(reg166) ?
                      $unsigned(reg77) : (~reg215))) ^~ $signed($unsigned((reg69 ^~ reg154)))) >= reg209);
            end
          reg226 <= $unsigned($signed((((&(8'hb3)) ? reg104 : (^~reg84)) ?
              ((reg56 ? reg224 : reg118) ?
                  (wire135 ?
                      (8'hb3) : reg198) : reg205[(3'h7):(3'h7)]) : $unsigned((8'haf)))));
          reg227 = {(8'hb8)};
          if ($unsigned($unsigned(({(~reg75), (reg142 >> reg109)} ?
              reg212[(4'hf):(4'hc)] : ($signed(forvar220) ? reg185 : reg217)))))
            begin
              reg228 <= $unsigned(reg203[(3'h5):(1'h1)]);
              reg229 <= (8'h9e);
              reg230 <= reg196[(4'h8):(1'h0)];
              reg231 = (7'h44);
            end
          else
            begin
              reg228 <= $signed(($unsigned($unsigned(((8'had) > reg166))) ?
                  (8'had) : reg107));
              reg231 = (reg229[(3'h5):(2'h3)] >>> $signed(reg69));
              reg232 = reg123[(4'h8):(2'h3)];
              reg233 <= reg225[(5'h10):(1'h1)];
            end
          if ($signed(reg208))
            begin
              reg234 <= $signed(wire40);
              reg235 = reg49[(2'h2):(1'h0)];
              reg236 <= $unsigned((8'hb6));
              reg237 = (^(8'h9c));
            end
          else
            begin
              reg235 = {reg128, reg204};
              reg237 = reg99[(1'h1):(1'h0)];
              reg238 = $unsigned((($signed((~|reg210)) ?
                  {$unsigned(reg186)} : $unsigned($unsigned((8'hb2)))) > ((^(forvar207 != reg228)) ?
                  ((reg74 ? reg225 : reg219) ?
                      (!reg225) : (reg93 ^~ reg211)) : (-reg55[(4'h8):(1'h1)]))));
              reg239 = $signed(($signed($signed(reg68[(1'h0):(1'h0)])) ?
                  (^reg93) : $unsigned(reg98)));
              reg240 <= $unsigned((|{$signed((reg84 ^~ reg154)),
                  reg213[(1'h1):(1'h0)]}));
            end
        end
      reg241 <= (^~(~&$signed((|$signed(reg206)))));
    end
  assign wire242 = reg142[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      reg243 <= (8'ha0);
      reg244 <= ({reg183,
          {reg192[(2'h2):(1'h1)],
              $unsigned(((8'ha7) < reg214))}} == ((((|reg99) + $signed(reg145)) == (-((8'hbc) | reg55))) ?
          (&(reg165[(2'h2):(1'h1)] ?
              reg228 : $unsigned(reg166))) : ($unsigned((~&(8'ha3))) <<< (^~reg216))));
      for (forvar245 = (1'h0); (forvar245 < (1'h0)); forvar245 = (forvar245 + (1'h1)))
        begin
          reg246 <= (|wire42[(4'hf):(4'hc)]);
          for (forvar247 = (1'h0); (forvar247 < (1'h0)); forvar247 = (forvar247 + (1'h1)))
            begin
              reg248 = reg215[(2'h3):(1'h0)];
              reg249 = $unsigned((|$unsigned(reg230[(4'h9):(3'h6)])));
              reg250 <= ((reg236 >= $signed($unsigned((^~reg133)))) * $unsigned($signed(wire38)));
              reg251 = $unsigned((reg146 ?
                  ($unsigned($unsigned(wire40)) & (8'ha9)) : (~$unsigned(reg85))));
              reg252 = $unsigned({($signed($signed(wire38)) ?
                      $unsigned((reg228 == (8'hb7))) : ((reg56 + reg186) ?
                          (reg192 - reg216) : (wire41 <<< reg192)))});
            end
        end
      reg253 = (((~^reg79) ~^ (reg175 ? reg139[(2'h2):(1'h1)] : reg211)) ?
          $signed((reg243[(5'h17):(5'h10)] ?
              $unsigned((!reg211)) : wire42)) : ((^~($signed(reg251) ?
                  reg214[(2'h2):(1'h1)] : $unsigned((8'h9f)))) ?
              (+((reg55 ? reg190 : reg196) ?
                  reg211[(1'h0):(1'h0)] : (~|reg77))) : $unsigned((reg80 ?
                  (reg208 ? reg145 : reg55) : $unsigned(reg90)))));
      for (forvar254 = (1'h0); (forvar254 < (3'h4)); forvar254 = (forvar254 + (1'h1)))
        begin
          reg255 <= $signed(reg128);
          reg256 = reg218;
          if ($signed(((($signed((8'ha8)) > reg234[(4'h9):(2'h3)]) ?
              reg178 : (wire38 ?
                  (reg203 ?
                      reg209 : reg104) : (reg68 > (8'hb6)))) >>> forvar254[(4'hf):(4'hc)])))
            begin
              reg257 <= (((~^$signed((reg240 ? reg142 : reg68))) ?
                      (reg117 ?
                          (7'h43) : (8'hb8)) : $unsigned($signed($signed(wire39)))) ?
                  ((^~reg110[(4'he):(4'hc)]) ?
                      reg146[(5'h14):(4'ha)] : {(^$signed(reg89)),
                          {(reg251 & reg153)}}) : reg223);
            end
          else
            begin
              reg257 <= reg198[(4'hb):(4'h8)];
              reg258 <= (|reg214[(2'h2):(1'h1)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg259 = reg52[(4'h9):(4'h9)];
    end
  always
    @(posedge clk) begin
      reg260 <= reg241;
      if (reg100[(1'h1):(1'h0)])
        begin
          reg261 <= (~&reg223);
          reg262 = ((~(+((reg243 ~^ reg209) || $signed((8'hae))))) ?
              (^reg79) : ($unsigned((((8'hab) || (7'h49)) ?
                  $unsigned(wire242) : reg96)) || $signed(wire39)));
        end
      else
        begin
          if ($signed(((reg262 >= {(reg46 ? reg223 : reg240),
              $signed(reg74)}) < (&($signed(reg222) ?
              (~^reg128) : (reg120 ? reg145 : reg146))))))
            begin
              reg262 = $unsigned(((reg133[(4'hf):(3'h7)] + (|$unsigned(reg68))) & $unsigned((~reg183[(2'h2):(1'h1)]))));
              reg263 = reg131[(4'h8):(3'h5)];
            end
          else
            begin
              reg262 = (reg192 ?
                  (&((reg243 == (8'ha6)) | {(reg74 ^~ reg100),
                      (reg216 ?
                          reg218 : reg96)})) : $signed($signed((+(reg261 ^ reg243)))));
              reg263 = $signed(((^(!$unsigned(reg205))) != reg46[(3'h4):(3'h4)]));
              reg264 <= (8'ha5);
              reg265 <= reg246;
            end
          for (forvar266 = (1'h0); (forvar266 < (1'h1)); forvar266 = (forvar266 + (1'h1)))
            begin
              reg267 <= (8'hbd);
            end
          reg268 <= reg145;
        end
      reg269 = $signed(((|(|$unsigned(reg104))) ?
          reg211[(4'hf):(1'h1)] : ({reg263[(3'h7):(3'h4)], (reg223 - reg126)} ?
              ((reg51 ? (8'h9d) : reg262) > {reg175}) : reg99[(3'h6):(2'h3)])));
      reg270 = (|(reg243 > reg258[(4'ha):(4'ha)]));
    end
  always
    @(posedge clk) begin
      if (reg261[(1'h0):(1'h0)])
        begin
          reg271 <= (wire140[(4'hb):(3'h4)] <<< (~({$signed(reg233)} & $signed((reg175 ?
              reg107 : reg203)))));
          reg272 <= $unsigned(($signed((reg175 > (reg171 ?
              reg172 : reg126))) == reg104[(3'h4):(1'h0)]));
          reg273 <= reg74[(3'h7):(1'h0)];
        end
      else
        begin
          for (forvar271 = (1'h0); (forvar271 < (2'h3)); forvar271 = (forvar271 + (1'h1)))
            begin
              reg272 <= (((~|wire41) ?
                      reg192 : $unsigned(($signed(reg51) >>> $unsigned(reg136)))) ?
                  ($signed(reg89[(3'h7):(1'h0)]) >>> (((reg156 <= wire140) ?
                          reg198 : (reg46 || (7'h40))) ?
                      {$signed(wire38), $signed(reg68)} : {$unsigned(reg211),
                          (reg224 | reg246)})) : reg169[(4'h9):(3'h6)]);
              reg274 = reg153;
              reg275 <= reg241[(5'h14):(1'h1)];
              reg276 <= (~|(^~$unsigned($unsigned((|reg236)))));
              reg277 <= $unsigned((reg276 ?
                  $unsigned(reg209) : (^$unsigned(reg226))));
            end
          reg278 <= ($signed(reg172) ~^ reg236);
        end
      reg279 = ({(~&($unsigned(reg128) >>> reg277))} < (!($signed(reg276[(5'h13):(4'hc)]) - $signed((reg233 ?
          (8'hab) : reg120)))));
    end
  always
    @(posedge clk) begin
      reg280 = $signed(($unsigned($unsigned(reg100[(3'h4):(1'h1)])) ?
          reg277 : (($signed(reg229) ? (~|reg72) : (8'hbe)) >> (~|((8'hb0) ?
              reg233 : reg77)))));
      reg281 = reg230[(4'ha):(1'h1)];
      if (($unsigned({reg89}) ?
          (reg211[(4'he):(4'hb)] | reg55) : reg202[(4'hb):(4'h8)]))
        begin
          reg282 <= {{reg267[(2'h3):(2'h3)], reg222},
              ($unsigned((^(reg215 != wire140))) * ((&reg142) ?
                  reg277 : $unsigned($signed(reg229))))};
          if (({reg202[(4'ha):(3'h5)]} ?
              (reg167[(3'h5):(1'h1)] ?
                  reg85[(4'hf):(4'hf)] : $unsigned((^~wire37))) : {((reg84[(1'h1):(1'h0)] ~^ (reg90 != (8'hbc))) << $unsigned($signed(reg145)))}))
            begin
              reg283 = (^~(~&$unsigned(((|reg136) ?
                  reg276 : reg156[(3'h4):(2'h2)]))));
              reg284 = ($signed(($signed(wire41) & (reg216[(4'h9):(3'h5)] ?
                  $unsigned(reg90) : $signed((8'ha0))))) ^ $signed(reg243));
              reg285 <= {$signed(reg190[(4'hf):(2'h3)])};
            end
          else
            begin
              reg283 = (^~$unsigned(reg272[(1'h1):(1'h0)]));
              reg285 <= {$unsigned(($signed($unsigned((7'h46))) != ((8'hb2) ?
                      reg142[(4'hc):(2'h2)] : reg84[(1'h0):(1'h0)]))),
                  {{{(reg278 ? reg264 : reg233)}}}};
              reg286 = ((reg167 >> (&wire38)) <<< reg84[(3'h5):(1'h0)]);
            end
          for (forvar287 = (1'h0); (forvar287 < (2'h3)); forvar287 = (forvar287 + (1'h1)))
            begin
              reg288 = wire41[(1'h0):(1'h0)];
            end
          reg289 = {reg218};
          reg290 = (reg178 ?
              reg214 : $unsigned({$unsigned(((8'hb6) || reg133))}));
        end
      else
        begin
          reg283 = reg55;
        end
    end
  assign wire291 = (({$unsigned((reg265 ? reg255 : wire39)),
                       (~{reg228, reg192})} || {$unsigned((reg99 ?
                           reg230 : reg203)),
                       reg178}) >= ((~wire41[(1'h0):(1'h0)]) ?
                       (8'hab) : reg75));
  always
    @(posedge clk) begin
      reg292 <= $signed((8'had));
      if ((((reg267 ~^ $unsigned(reg107)) ?
          $unsigned({$unsigned((7'h45)),
              (-reg185)}) : ({(reg258 >> (8'hac))} << (+{reg192}))) + $signed(reg120[(1'h0):(1'h0)])))
        begin
          if ((reg202 && (($unsigned(reg133[(4'hd):(1'h1)]) ?
                  $unsigned((reg276 ?
                      reg84 : (8'ha0))) : (reg136[(3'h6):(1'h1)] ?
                      (|reg169) : reg260)) ?
              $signed($signed($signed(wire39))) : (($signed(reg98) ?
                      wire140[(4'h9):(4'h8)] : {(8'ha8), reg292}) ?
                  $signed(wire291) : reg255[(3'h7):(3'h6)]))))
            begin
              reg293 <= (((8'hac) ?
                  reg68 : $unsigned($signed(wire41[(1'h0):(1'h0)]))) << reg273[(3'h4):(1'h0)]);
              reg294 <= reg69[(1'h1):(1'h0)];
              reg295 = ($unsigned(reg226) ?
                  $unsigned({$unsigned(((7'h41) ? (8'hb3) : (8'had))),
                      (8'hac)}) : (+($signed({wire158, (8'hbf)}) ?
                      $unsigned(wire291) : $signed(reg219[(1'h1):(1'h0)]))));
              reg296 = wire42;
              reg297 = ($unsigned(($signed(reg123) ?
                  reg93[(1'h0):(1'h0)] : (!(7'h49)))) < reg294);
            end
          else
            begin
              reg295 = (8'ha1);
            end
          for (forvar298 = (1'h0); (forvar298 < (1'h1)); forvar298 = (forvar298 + (1'h1)))
            begin
              reg299 = (reg192[(3'h4):(3'h4)] == ($unsigned(($signed((8'hb0)) ?
                  $unsigned(reg93) : (reg222 ^ reg46))) || {$signed(reg275[(2'h2):(2'h2)])}));
              reg300 = (&$unsigned(($unsigned(reg153[(3'h4):(1'h0)]) ?
                  (~$signed(reg139)) : reg261)));
              reg301 <= {reg169};
              reg302 <= {reg166};
            end
          reg303 = reg136;
          for (forvar304 = (1'h0); (forvar304 < (1'h1)); forvar304 = (forvar304 + (1'h1)))
            begin
              reg305 <= (($unsigned(reg56) <= (reg133 ?
                  reg85 : reg302)) >> wire38[(4'h9):(3'h6)]);
            end
        end
      else
        begin
          reg293 <= wire40[(1'h0):(1'h0)];
          if ($unsigned($unsigned(reg136)))
            begin
              reg294 <= $signed((~^$unsigned((~|(~&reg302)))));
            end
          else
            begin
              reg294 <= ({(-(8'h9f)),
                      ({$signed(reg267)} + (!(reg185 << (8'hb1))))} ?
                  $unsigned(((^~reg136[(3'h7):(2'h3)]) ?
                      reg257 : $unsigned($signed(reg215)))) : reg84);
              reg295 = reg223[(3'h7):(3'h6)];
              reg296 = $signed((({$unsigned(reg117), {reg276}} ?
                      reg77[(3'h5):(3'h5)] : reg198[(4'he):(3'h4)]) ?
                  $unsigned($signed(((8'had) ?
                      reg46 : wire140))) : reg51[(1'h0):(1'h0)]));
              reg297 = reg46[(1'h0):(1'h0)];
              reg298 <= {reg216};
            end
        end
    end
  always
    @(posedge clk) begin
      reg306 <= (~&$unsigned(reg292));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module947  (y, clk, wire951, wire950, wire949, wire948);
  output wire [(32'hc2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire951;
  input wire [(4'hf):(1'h0)] wire950;
  input wire signed [(4'h8):(1'h0)] wire949;
  input wire [(4'h9):(1'h0)] wire948;
  wire signed [(3'h5):(1'h0)] wire964;
  wire [(5'h13):(1'h0)] wire963;
  wire signed [(4'he):(1'h0)] wire955;
  wire signed [(4'hc):(1'h0)] wire954;
  wire [(5'h14):(1'h0)] wire953;
  wire [(5'h12):(1'h0)] wire952;
  reg signed [(3'h4):(1'h0)] reg961 = (1'h0);
  reg [(4'hc):(1'h0)] reg960 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg957 = (1'h0);
  reg [(5'h10):(1'h0)] reg956 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg962 = (1'h0);
  reg [(5'h14):(1'h0)] reg959 = (1'h0);
  reg [(5'h17):(1'h0)] reg958 = (1'h0);
  assign y = {wire964,
                 wire963,
                 wire955,
                 wire954,
                 wire953,
                 wire952,
                 reg961,
                 reg960,
                 reg957,
                 reg956,
                 reg962,
                 reg959,
                 reg958,
                 (1'h0)};
  assign wire952 = $signed(wire950);
  assign wire953 = $unsigned(wire949);
  assign wire954 = {($signed((wire953 ?
                           $unsigned(wire953) : wire949)) && (wire948[(2'h2):(2'h2)] ?
                           wire949[(3'h5):(2'h2)] : $unsigned($signed(wire948)))),
                       wire950[(4'hb):(3'h5)]};
  assign wire955 = $signed({$unsigned($signed((wire954 ^ wire948))),
                       (wire950 ^ (~^wire953[(3'h6):(2'h2)]))});
  always
    @(posedge clk) begin
      reg956 <= ($unsigned($unsigned((wire950 ?
          (~|wire950) : (wire948 ?
              wire951 : wire949)))) <= ($signed(wire951[(4'ha):(1'h0)]) ?
          $signed(((wire954 ?
              wire955 : wire955) == wire955[(3'h6):(3'h5)])) : wire953));
      reg957 <= ($unsigned(wire953[(5'h10):(4'hf)]) ?
          $unsigned(wire953) : $signed($unsigned(wire952[(4'hc):(1'h0)])));
      reg958 = (($unsigned((wire948 >= (reg957 >= reg956))) + ({(|(8'hae)),
              (wire953 ? wire951 : reg957)} ?
          ({wire951, wire949} ?
              {wire949, wire950} : {wire949, reg956}) : {(reg956 - wire949),
              ((8'h9d) ~^ wire948)})) >>> (~|{$unsigned(wire955[(3'h5):(1'h1)])}));
      reg959 = (+(^~wire950[(4'hb):(4'ha)]));
    end
  always
    @(posedge clk) begin
      reg960 <= $unsigned(((~|$unsigned((wire948 ?
          (8'hb5) : (8'ha4)))) | wire952[(5'h11):(5'h11)]));
      reg961 <= (wire952 ?
          reg957[(4'hb):(3'h7)] : ($signed(((wire952 ~^ (7'h49)) || $signed(reg956))) >= wire948));
      reg962 = reg961;
    end
  assign wire963 = (($signed(((wire949 ?
                           wire955 : wire949) >= reg956[(4'he):(3'h6)])) == reg961[(2'h2):(1'h1)]) ?
                       $unsigned(reg957[(2'h2):(1'h1)]) : (($signed(reg960[(2'h2):(1'h1)]) || reg956[(4'h8):(3'h7)]) <= wire953[(4'h8):(3'h7)]));
  assign wire964 = {reg961};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module533
#(parameter param914 = (((({(8'hbf)} ? ((8'hbe) != (8'h9e)) : ((8'ha4) ? (7'h43) : (8'ha5))) >>> {((8'hab) & (8'hbd))}) ? ((((8'hab) && (7'h44)) ^~ ((8'ha9) > (8'ha5))) ? (((8'h9d) < (7'h47)) < (^(7'h43))) : (~^((8'hb6) != (8'hbf)))) : ((&((8'ha7) ? (8'hbc) : (8'hba))) ? {((8'haa) >> (8'had))} : (~&((8'hb7) ? (8'hb7) : (7'h46))))) - (((((8'h9e) ? (8'hbf) : (8'hac)) ? (^(8'hb7)) : {(8'ha1), (7'h42)}) && ((7'h43) ^~ (^(8'had)))) | (~^(~&(-(8'ha7)))))))
(y, clk, wire534, wire535, wire536, wire537);
  output wire [(32'h646):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h16):(1'h0)] wire534;
  input wire signed [(4'hd):(1'h0)] wire535;
  input wire signed [(5'h16):(1'h0)] wire536;
  input wire [(2'h3):(1'h0)] wire537;
  wire [(3'h7):(1'h0)] wire913;
  wire signed [(4'hb):(1'h0)] wire911;
  wire [(4'hd):(1'h0)] wire910;
  wire signed [(4'hc):(1'h0)] wire738;
  wire [(5'h18):(1'h0)] wire740;
  wire signed [(4'hf):(1'h0)] wire759;
  wire signed [(5'h12):(1'h0)] wire760;
  wire signed [(3'h7):(1'h0)] wire778;
  wire signed [(5'h13):(1'h0)] wire794;
  wire [(5'h17):(1'h0)] wire801;
  wire [(3'h4):(1'h0)] wire802;
  wire [(2'h2):(1'h0)] wire908;
  reg signed [(5'h11):(1'h0)] reg912 = (1'h0);
  reg [(5'h14):(1'h0)] reg577 = (1'h0);
  reg [(5'h11):(1'h0)] reg576 = (1'h0);
  reg [(5'h10):(1'h0)] reg575 = (1'h0);
  reg [(5'h11):(1'h0)] reg574 = (1'h0);
  reg [(5'h11):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg568 = (1'h0);
  reg [(3'h4):(1'h0)] reg567 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg566 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg563 = (1'h0);
  reg [(5'h14):(1'h0)] reg561 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg560 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg558 = (1'h0);
  reg [(3'h7):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg554 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg545 = (1'h0);
  reg [(3'h7):(1'h0)] reg544 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg542 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg539 = (1'h0);
  reg [(5'h17):(1'h0)] reg538 = (1'h0);
  reg [(5'h11):(1'h0)] reg743 = (1'h0);
  reg [(2'h3):(1'h0)] reg745 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg750 = (1'h0);
  reg [(2'h3):(1'h0)] reg752 = (1'h0);
  reg [(5'h15):(1'h0)] reg753 = (1'h0);
  reg [(4'h9):(1'h0)] reg754 = (1'h0);
  reg [(4'ha):(1'h0)] reg751 = (1'h0);
  reg [(5'h18):(1'h0)] reg757 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg761 = (1'h0);
  reg [(3'h7):(1'h0)] reg766 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg767 = (1'h0);
  reg [(4'hc):(1'h0)] reg769 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg770 = (1'h0);
  reg [(5'h16):(1'h0)] reg772 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg765 = (1'h0);
  reg [(5'h11):(1'h0)] reg771 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg774 = (1'h0);
  reg [(3'h4):(1'h0)] reg775 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg776 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg777 = (1'h0);
  reg [(4'hc):(1'h0)] reg783 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg784 = (1'h0);
  reg [(3'h4):(1'h0)] reg785 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg789 = (1'h0);
  reg [(4'he):(1'h0)] reg790 = (1'h0);
  reg [(4'hf):(1'h0)] reg792 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg799 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg800 = (1'h0);
  reg [(5'h16):(1'h0)] reg803 = (1'h0);
  reg [(5'h15):(1'h0)] reg798 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg797 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar796 = (1'h0);
  reg [(3'h6):(1'h0)] reg795 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg793 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg791 = (1'h0);
  reg [(5'h15):(1'h0)] reg788 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg787 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg786 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg782 = (1'h0);
  reg [(4'hc):(1'h0)] reg781 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg780 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar779 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg773 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg763 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar771 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg768 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar765 = (1'h0);
  reg [(3'h7):(1'h0)] reg764 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar763 = (1'h0);
  reg signed [(4'he):(1'h0)] reg762 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg758 = (1'h0);
  reg [(4'ha):(1'h0)] reg756 = (1'h0);
  reg [(3'h6):(1'h0)] reg755 = (1'h0);
  reg [(5'h15):(1'h0)] forvar751 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg749 = (1'h0);
  reg [(5'h13):(1'h0)] reg748 = (1'h0);
  reg [(5'h17):(1'h0)] forvar747 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg746 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar744 = (1'h0);
  reg [(4'hc):(1'h0)] forvar742 = (1'h0);
  reg [(5'h18):(1'h0)] reg741 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg573 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg572 = (1'h0);
  reg [(5'h10):(1'h0)] reg571 = (1'h0);
  reg [(3'h4):(1'h0)] reg569 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg565 = (1'h0);
  reg [(5'h13):(1'h0)] forvar564 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg562 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar559 = (1'h0);
  reg [(4'ha):(1'h0)] reg557 = (1'h0);
  reg [(4'h9):(1'h0)] reg555 = (1'h0);
  reg [(2'h3):(1'h0)] reg553 = (1'h0);
  reg [(4'hc):(1'h0)] forvar552 = (1'h0);
  reg [(5'h18):(1'h0)] reg551 = (1'h0);
  reg [(5'h11):(1'h0)] reg550 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg549 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg548 = (1'h0);
  reg [(2'h3):(1'h0)] reg547 = (1'h0);
  reg [(5'h13):(1'h0)] forvar546 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg543 = (1'h0);
  reg [(3'h7):(1'h0)] reg541 = (1'h0);
  reg signed [(4'he):(1'h0)] reg540 = (1'h0);
  assign y = {wire913,
                 wire911,
                 wire910,
                 wire738,
                 wire740,
                 wire759,
                 wire760,
                 wire778,
                 wire794,
                 wire801,
                 wire802,
                 wire908,
                 reg912,
                 reg577,
                 reg576,
                 reg575,
                 reg574,
                 reg570,
                 reg568,
                 reg567,
                 reg566,
                 reg563,
                 reg561,
                 reg560,
                 reg558,
                 reg556,
                 reg554,
                 reg545,
                 reg544,
                 reg542,
                 reg539,
                 reg538,
                 reg743,
                 reg745,
                 reg750,
                 reg752,
                 reg753,
                 reg754,
                 reg751,
                 reg757,
                 reg761,
                 reg766,
                 reg767,
                 reg769,
                 reg770,
                 reg772,
                 reg765,
                 reg771,
                 reg774,
                 reg775,
                 reg776,
                 reg777,
                 reg783,
                 reg784,
                 reg785,
                 reg789,
                 reg790,
                 reg792,
                 reg799,
                 reg800,
                 reg803,
                 reg798,
                 reg797,
                 forvar796,
                 reg795,
                 reg793,
                 reg791,
                 reg788,
                 reg787,
                 reg786,
                 reg782,
                 reg781,
                 reg780,
                 forvar779,
                 reg773,
                 reg763,
                 forvar771,
                 reg768,
                 forvar765,
                 reg764,
                 forvar763,
                 reg762,
                 reg758,
                 reg756,
                 reg755,
                 forvar751,
                 reg749,
                 reg748,
                 forvar747,
                 reg746,
                 forvar744,
                 forvar742,
                 reg741,
                 reg573,
                 reg572,
                 reg571,
                 reg569,
                 reg565,
                 forvar564,
                 reg562,
                 forvar559,
                 reg557,
                 reg555,
                 reg553,
                 forvar552,
                 reg551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 forvar546,
                 reg543,
                 reg541,
                 reg540,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg538 <= wire534;
      reg539 <= {((wire535 ^ wire536[(4'h8):(2'h3)]) == (wire535[(1'h1):(1'h1)] >>> ((8'hbb) == $signed(reg538)))),
          ((^(|$unsigned((7'h43)))) || $signed(($unsigned(wire536) ?
              {wire534} : (7'h44))))};
      if (wire534)
        begin
          reg540 = $signed({wire535});
        end
      else
        begin
          reg540 = $unsigned($unsigned((wire536 ?
              ((wire535 * reg538) <= (wire535 | wire537)) : ((wire534 + wire535) * wire535))));
          if (((wire535 && reg538) || ($signed(wire537) ? {(8'hb8)} : (7'h4a))))
            begin
              reg541 = $signed((~^reg540[(3'h6):(2'h2)]));
            end
          else
            begin
              reg541 = {(-((^(reg541 ? wire536 : wire537)) ?
                      ($unsigned(reg538) << (reg540 <= reg539)) : (~|reg540[(3'h7):(1'h1)]))),
                  reg541[(1'h1):(1'h0)]};
              reg542 <= (reg541[(3'h6):(1'h0)] ?
                  (+(wire534 ?
                      $unsigned(reg540) : $signed($signed(reg541)))) : $signed((+(reg539[(3'h5):(1'h0)] || $signed(reg541)))));
              reg543 = $signed(reg542);
              reg544 <= $signed(({($unsigned(reg543) ^~ reg541[(2'h3):(2'h2)]),
                      reg539[(4'ha):(2'h2)]} ?
                  (((wire534 << reg540) <= (7'h49)) ?
                      {((8'h9f) ?
                              reg543 : (8'hb0))} : wire535[(4'h9):(3'h7)]) : $unsigned(wire537)));
              reg545 <= $signed(wire534);
            end
          for (forvar546 = (1'h0); (forvar546 < (3'h4)); forvar546 = (forvar546 + (1'h1)))
            begin
              reg547 = (!$signed(((7'h44) ? wire537 : (!{wire534, reg539}))));
              reg548 = reg541;
              reg549 = (~(~{($signed(reg545) | reg543), reg543}));
              reg550 = {$signed({$signed((reg543 ? reg539 : reg541))}),
                  ((|$signed(wire534[(4'ha):(3'h4)])) ^~ ($signed(forvar546) ?
                      reg540[(4'ha):(4'h8)] : (~^((8'hb6) ?
                          reg544 : reg538))))};
              reg551 = reg543;
            end
          for (forvar552 = (1'h0); (forvar552 < (1'h0)); forvar552 = (forvar552 + (1'h1)))
            begin
              reg553 = wire537;
              reg554 <= ({$unsigned(($signed(reg543) ?
                      (~^forvar546) : $unsigned(reg540))),
                  reg551} ^~ (reg548 <<< $signed(forvar546)));
              reg555 = (($unsigned((forvar552 ?
                  (wire534 & reg549) : $unsigned(reg554))) < reg544) & forvar552[(1'h0):(1'h0)]);
              reg556 <= {(^~reg540[(3'h5):(3'h5)])};
              reg557 = (~^reg550[(3'h4):(1'h0)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg558 <= $unsigned($signed(reg544));
      for (forvar559 = (1'h0); (forvar559 < (2'h3)); forvar559 = (forvar559 + (1'h1)))
        begin
          reg560 <= $unsigned(((+($unsigned(reg538) ?
                  (~|reg545) : (~(8'ha2)))) ?
              $signed(reg538[(2'h2):(2'h2)]) : ((^{reg544}) ?
                  ((reg545 <= (7'h42)) > (reg545 ?
                      reg545 : reg544)) : ((wire537 ? (8'hbd) : reg545) ?
                      $signed(reg544) : (reg538 + wire534)))));
          reg561 <= reg538[(5'h14):(5'h11)];
          reg562 = $signed(((~^(|((8'hbe) * (7'h4a)))) && $signed((~^$signed(wire536)))));
        end
      reg563 <= wire535[(3'h5):(3'h4)];
      for (forvar564 = (1'h0); (forvar564 < (3'h4)); forvar564 = (forvar564 + (1'h1)))
        begin
          if (forvar564[(3'h7):(3'h5)])
            begin
              reg565 = (~|((~&reg561[(5'h14):(5'h10)]) | reg556[(2'h3):(1'h0)]));
              reg566 <= $unsigned(wire535[(4'hb):(4'ha)]);
              reg567 <= $signed((((reg544 * {wire536, reg565}) ?
                      wire535[(4'ha):(1'h0)] : $signed((reg544 ?
                          reg563 : reg561))) ?
                  {($unsigned(forvar559) ?
                          wire535 : $unsigned((8'hb1)))} : reg538[(3'h6):(3'h4)]));
            end
          else
            begin
              reg566 <= reg566[(2'h2):(1'h1)];
            end
          if ((((~&($unsigned(reg542) ?
              (-reg539) : wire537)) >= ((forvar559[(2'h2):(1'h0)] ?
              $signed(forvar564) : $signed(reg562)) & (reg558[(1'h1):(1'h1)] ?
              $unsigned(reg539) : (~^reg565)))) | ($unsigned(wire537) ?
              (reg542 >>> reg566) : (8'haf))))
            begin
              reg568 <= {reg563[(4'hb):(3'h5)]};
            end
          else
            begin
              reg569 = $unsigned((^~(~&$signed($unsigned(reg544)))));
              reg570 <= reg568;
              reg571 = $unsigned($signed(($unsigned((^~reg569)) ?
                  (8'hab) : $unsigned($unsigned(reg569)))));
              reg572 = $unsigned($unsigned((($unsigned(reg560) - ((8'ha2) > forvar559)) > ((wire537 ?
                      wire537 : wire534) ?
                  reg567[(1'h1):(1'h1)] : {(8'hae), reg566}))));
            end
          reg573 = $signed((reg554 ^~ ($unsigned($signed((8'hac))) && ((reg554 ?
              (8'hbe) : reg567) <= (reg542 ? (8'hb4) : wire534)))));
          if (($signed(((|$unsigned(reg558)) && $signed((|reg567)))) ?
              (((&(~^forvar564)) ?
                  (7'h44) : reg562[(4'ha):(3'h7)]) * (!($unsigned(reg554) ?
                  $unsigned(reg565) : (reg554 ?
                      reg538 : reg539)))) : ($unsigned(($signed((8'hb6)) ?
                  (-reg560) : $signed(reg566))) >>> reg573[(1'h1):(1'h1)])))
            begin
              reg574 <= $unsigned($unsigned({({reg561, reg538} ?
                      (~^reg538) : (^(7'h48)))}));
            end
          else
            begin
              reg574 <= reg545[(3'h7):(3'h6)];
              reg575 <= wire537;
              reg576 <= (~|$unsigned($unsigned((reg568 - $unsigned(reg573)))));
              reg577 <= reg565[(4'hc):(3'h4)];
            end
        end
    end
  module578 #() modinst739 (.wire582(reg542), .y(wire738), .wire583(reg574), .wire581(wire534), .clk(clk), .wire580(reg558), .wire579(wire536));
  assign wire740 = $signed(reg570);
  always
    @(posedge clk) begin
      reg741 = ((reg567[(2'h2):(1'h0)] ?
              (reg554[(5'h13):(3'h4)] || reg576) : (8'h9e)) ?
          $signed(reg570[(4'hf):(4'h8)]) : (&$signed((+reg556))));
      for (forvar742 = (1'h0); (forvar742 < (3'h4)); forvar742 = (forvar742 + (1'h1)))
        begin
          reg743 <= reg554;
        end
      for (forvar744 = (1'h0); (forvar744 < (1'h0)); forvar744 = (forvar744 + (1'h1)))
        begin
          reg745 <= {(((~|$unsigned(reg542)) ?
                  $unsigned((reg575 || reg743)) : $signed((8'hbe))) ^~ ($signed(reg561[(3'h5):(2'h2)]) ?
                  wire740 : $signed($unsigned(reg576)))),
              (reg561[(5'h10):(4'hd)] < (&{reg558[(2'h3):(2'h2)]}))};
          reg746 = $signed($unsigned((reg539[(3'h6):(1'h0)] ?
              (~|(-(8'ha5))) : $unsigned(reg566[(4'ha):(3'h6)]))));
          for (forvar747 = (1'h0); (forvar747 < (1'h1)); forvar747 = (forvar747 + (1'h1)))
            begin
              reg748 = {(7'h40)};
              reg749 = $unsigned(reg538);
            end
        end
    end
  always
    @(posedge clk) begin
      reg750 <= $unsigned((($unsigned(reg542) ?
              (reg566[(2'h3):(1'h1)] ?
                  (+(8'ha3)) : $signed(wire536)) : {(^~reg558)}) ?
          wire537 : $unsigned({$signed(reg577)})));
      if ($signed(reg560[(3'h4):(1'h0)]))
        begin
          for (forvar751 = (1'h0); (forvar751 < (1'h1)); forvar751 = (forvar751 + (1'h1)))
            begin
              reg752 <= (^wire537[(1'h0):(1'h0)]);
              reg753 <= reg750;
              reg754 <= ($signed($signed(reg574[(5'h11):(1'h1)])) ?
                  reg539 : {reg577});
            end
          reg755 = wire738[(4'h9):(4'h8)];
        end
      else
        begin
          if ($signed($unsigned({reg560[(4'he):(4'h8)]})))
            begin
              reg751 <= reg754;
              reg752 <= ($signed($unsigned({((7'h47) ? (8'h9f) : (8'h9c)),
                      (~^reg752)})) ?
                  $unsigned({reg755[(1'h1):(1'h1)],
                      reg558}) : ((($signed(reg566) != ((7'h43) ?
                      wire738 : reg538)) > reg753[(5'h15):(1'h0)]) || reg570));
            end
          else
            begin
              reg751 <= ((~|reg566[(3'h4):(3'h4)]) <<< (reg568 ?
                  $signed(((reg566 ? reg561 : (8'haf)) ?
                      $unsigned(reg576) : (forvar751 ?
                          reg538 : reg539))) : ($unsigned((wire537 + (8'ha9))) > (((7'h45) || reg566) ?
                      (~wire740) : (+reg575)))));
            end
        end
      reg756 = reg753[(5'h13):(3'h4)];
      reg757 <= ((+(reg561 >= ((+wire740) ?
          $unsigned(reg542) : (reg574 && reg575)))) << (({reg538[(4'he):(4'he)]} ^ (8'hb7)) ^~ reg567));
      reg758 = reg754;
    end
  assign wire759 = reg556[(3'h5):(3'h5)];
  assign wire760 = (reg757[(4'hd):(4'hb)] > {(8'hac), reg558});
  always
    @(posedge clk) begin
      if ($signed($signed((~(&{(8'ha9)})))))
        begin
          if ($signed(((8'h9e) | (8'haf))))
            begin
              reg761 <= reg751;
              reg762 = $signed($signed(($signed(reg577) << $signed(reg560[(4'hf):(3'h7)]))));
            end
          else
            begin
              reg762 = reg554;
            end
          for (forvar763 = (1'h0); (forvar763 < (1'h1)); forvar763 = (forvar763 + (1'h1)))
            begin
              reg764 = $unsigned($signed($unsigned(wire759)));
            end
          for (forvar765 = (1'h0); (forvar765 < (2'h2)); forvar765 = (forvar765 + (1'h1)))
            begin
              reg766 <= $unsigned(wire535);
              reg767 <= ((8'hb6) ?
                  $signed({(((8'h9c) ? reg567 : (8'hbd)) ?
                          (~|reg745) : $unsigned(wire536)),
                      $unsigned($signed(wire535))}) : $unsigned((wire759[(4'ha):(4'h9)] ?
                      ({reg577} ?
                          $unsigned(reg538) : wire534[(4'ha):(2'h2)]) : $unsigned((reg545 ?
                          reg576 : reg561)))));
              reg768 = reg560;
              reg769 <= reg577[(4'h9):(4'h9)];
              reg770 <= reg556[(2'h3):(1'h0)];
            end
          for (forvar771 = (1'h0); (forvar771 < (2'h3)); forvar771 = (forvar771 + (1'h1)))
            begin
              reg772 <= {reg570[(3'h6):(2'h3)]};
            end
        end
      else
        begin
          if ({reg574})
            begin
              reg762 = reg574[(2'h2):(1'h0)];
              reg763 = (8'hae);
              reg765 <= ((reg561 ?
                      (reg576 < $unsigned(reg576[(4'h9):(3'h7)])) : {reg761}) ?
                  ((reg563 ? reg576 : (~&reg769[(2'h3):(1'h1)])) ?
                      {(reg750 ? (reg751 > (8'hb6)) : (~&(7'h45))),
                          wire537} : ({(forvar763 + reg757),
                          $unsigned(reg574)} == (&(^~(8'hbb))))) : reg556[(1'h0):(1'h0)]);
              reg768 = $unsigned($signed((^{{reg566, reg765},
                  (wire740 ? (8'hb3) : reg762)})));
            end
          else
            begin
              reg762 = reg556;
              reg763 = $signed(({{$signed(reg554), reg751},
                      ({forvar763, reg751} ? $signed((7'h4a)) : (8'hb3))} ?
                  {((reg768 ? (8'hb1) : reg772) - ((8'hbb) ?
                          reg561 : reg566))} : ((((8'ha5) ? wire535 : reg538) ?
                          {reg576, reg752} : reg577) ?
                      ($signed(forvar771) ?
                          $signed(reg768) : {reg767,
                              reg566}) : (reg743[(4'h9):(3'h5)] ?
                          ((8'hba) >= forvar771) : reg538))));
            end
          if ((&$signed($unsigned({{(8'ha8)}, (~&forvar763)}))))
            begin
              reg769 <= ($unsigned($unsigned(reg568[(4'he):(4'he)])) || {reg766[(2'h3):(2'h3)]});
              reg770 <= $unsigned(reg545);
              reg771 <= {$signed(wire738)};
              reg773 = $signed($signed((((!reg577) ^ {reg766, (7'h40)}) ?
                  reg745[(1'h0):(1'h0)] : (((8'hbd) < (8'ha5)) + (reg768 ?
                      reg752 : reg558)))));
            end
          else
            begin
              reg769 <= (~^(((reg568 > (reg563 ?
                      reg574 : reg560)) && (((8'ha1) ?
                      reg751 : reg574) <<< $unsigned((8'hb7)))) ?
                  (+($unsigned(wire534) != (reg770 >>> reg567))) : $signed(((forvar765 & reg556) <<< (wire759 ?
                      reg750 : forvar763)))));
              reg770 <= (reg570[(2'h3):(2'h3)] ?
                  wire740 : {{$signed($unsigned(reg772))},
                      {((~&(7'h41)) >>> {reg539, reg570})}});
              reg773 = (($unsigned(reg752) && $unsigned($signed(reg544[(1'h1):(1'h1)]))) ?
                  reg561[(2'h3):(2'h3)] : $signed(forvar771));
            end
        end
    end
  always
    @(posedge clk) begin
      reg774 <= {((((!reg770) ?
                  reg577[(4'hf):(4'hb)] : (wire740 ?
                      reg570 : wire760)) <= $unsigned((reg570 ?
                  reg542 : reg769))) ?
              reg563 : $signed((~^(8'hb7)))),
          ({$unsigned((reg772 ? reg754 : reg558)),
                  {(wire536 >> reg769), {(8'h9f)}}} ?
              $unsigned((+reg576)) : $signed(($signed(wire760) ?
                  reg568[(4'ha):(3'h4)] : reg554)))};
      reg775 <= wire534[(5'h10):(4'hd)];
      reg776 <= reg766[(1'h1):(1'h0)];
      reg777 <= (((~|((^reg771) ~^ {wire759})) ?
          {((&reg539) ?
                  {wire534} : reg545[(2'h3):(2'h2)])} : ({$signed(wire534),
                  wire537} ?
              $unsigned(reg766[(2'h3):(1'h1)]) : ((reg561 ? reg558 : wire740) ?
                  (wire535 << (8'hb7)) : $signed(reg766)))) ^~ wire738[(3'h5):(1'h0)]);
    end
  assign wire778 = ((!reg775[(2'h2):(1'h0)]) ?
                       reg563[(1'h1):(1'h1)] : wire537[(1'h1):(1'h1)]);
  always
    @(posedge clk) begin
      for (forvar779 = (1'h0); (forvar779 < (1'h1)); forvar779 = (forvar779 + (1'h1)))
        begin
          if ((8'hb0))
            begin
              reg780 = ({(~&reg570[(5'h10):(1'h0)])} ?
                  $unsigned((((|(8'hb7)) * $signed((8'hb0))) ^ $signed((reg767 || reg751)))) : (((&(|(8'hb2))) || (^reg542)) ^ reg568[(4'hc):(3'h5)]));
              reg781 = {wire738[(4'h9):(4'h9)], (~reg750[(1'h1):(1'h1)])};
              reg782 = {(^~reg753)};
            end
          else
            begin
              reg780 = ($unsigned((|{{reg781, reg576},
                  reg776[(3'h4):(3'h4)]})) + (wire738[(2'h2):(1'h0)] ?
                  $signed($unsigned((reg567 ?
                      reg576 : reg752))) : ($unsigned($unsigned(reg757)) - wire738[(4'hb):(4'h8)])));
              reg783 <= reg568;
              reg784 <= (-$signed($signed(((reg777 ? reg757 : reg561) ?
                  ((8'h9e) & reg575) : (reg757 + reg542)))));
            end
          reg785 <= (~$unsigned({((reg752 ? reg784 : reg750) >= (wire760 ?
                  reg568 : reg558)),
              ((+(8'hbb)) & ((8'ha3) ? reg765 : reg761))}));
          reg786 = $unsigned(wire778[(1'h1):(1'h0)]);
          reg787 = ((reg776[(3'h5):(2'h3)] != reg775) <= $signed(reg751[(3'h4):(2'h2)]));
          if ($unsigned($unsigned(reg560[(4'hd):(4'h9)])))
            begin
              reg788 = (reg783 + reg781);
              reg789 <= {(^~(+({(8'ha1)} + (8'h9c))))};
              reg790 <= (^reg765);
              reg791 = (((^~$signed((reg776 ?
                  reg568 : wire535))) > $signed($unsigned(reg783))) ^ (reg753 ?
                  (^~reg558) : reg750));
              reg792 <= (-(|$signed($signed(reg568[(1'h1):(1'h1)]))));
            end
          else
            begin
              reg789 <= (((((wire778 <<< reg570) & wire760) >> $signed((~&reg566))) ?
                  $signed(($signed(reg750) ?
                      (|reg783) : $unsigned((8'h9d)))) : reg563[(4'hb):(1'h1)]) && (reg575[(4'hb):(4'hb)] ?
                  wire778 : reg753[(5'h15):(3'h7)]));
              reg791 = (~|reg772);
              reg792 <= ({$unsigned(reg563)} <= (7'h49));
              reg793 = {(reg770[(2'h3):(1'h1)] & ($unsigned((reg781 ?
                          reg766 : reg766)) ?
                      reg538 : (~|$unsigned((8'h9e))))),
                  (^$unsigned((7'h41)))};
            end
        end
    end
  assign wire794 = $unsigned((reg777[(3'h6):(3'h5)] ^~ wire759[(3'h5):(3'h4)]));
  always
    @(posedge clk) begin
      reg795 = $unsigned($signed((wire740 || reg769)));
      for (forvar796 = (1'h0); (forvar796 < (1'h0)); forvar796 = (forvar796 + (1'h1)))
        begin
          if (((reg771[(1'h0):(1'h0)] ?
                  (((|reg770) & $unsigned(reg775)) | $signed(wire760[(4'hc):(4'ha)])) : $unsigned(reg790)) ?
              $signed((~^$signed((forvar796 <= (8'hae))))) : (~^(~$signed(reg753)))))
            begin
              reg797 = (reg554[(5'h14):(2'h2)] * $unsigned($unsigned((reg769[(4'ha):(4'h9)] ?
                  (reg767 ? reg754 : reg751) : reg784[(2'h2):(2'h2)]))));
              reg798 = $signed((reg542 <<< {reg743, forvar796[(2'h3):(2'h2)]}));
              reg799 <= ($signed((wire740 ?
                  (~^(reg577 ?
                      (8'haa) : reg798)) : ((reg777 <<< wire534) << wire536[(4'he):(4'he)]))) <= $unsigned($signed($signed(reg570[(2'h2):(1'h0)]))));
            end
          else
            begin
              reg799 <= $signed(reg577[(3'h5):(2'h3)]);
            end
          reg800 <= ($unsigned($signed(reg783)) ^~ ($unsigned({$unsigned(reg539)}) ?
              (|reg568[(3'h5):(1'h1)]) : $unsigned($unsigned($unsigned(reg792)))));
        end
    end
  assign wire801 = (((7'h40) ?
                       $signed({(reg576 ? wire534 : (7'h43)),
                           $signed(reg750)}) : {(reg800 - reg568)}) + wire778[(1'h0):(1'h0)]);
  assign wire802 = $unsigned($signed((wire537 != {$unsigned(reg556),
                       $unsigned(wire759)})));
  always
    @(posedge clk) begin
      reg803 <= ($signed($unsigned((reg568[(4'hf):(4'h8)] > ((8'h9d) ?
          reg561 : reg754)))) >>> $signed($signed($unsigned(((8'haf) ?
          reg777 : reg800)))));
    end
  module804 #() modinst909 (.wire807(wire738), .wire805(wire778), .wire806(reg771), .clk(clk), .y(wire908), .wire808(wire801));
  assign wire910 = reg544[(3'h4):(2'h3)];
  assign wire911 = {$unsigned(($signed((reg785 ?
                           wire738 : wire759)) & reg771))};
  always
    @(posedge clk) begin
      reg912 <= reg767;
    end
  assign wire913 = reg556[(2'h2):(1'h1)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module804  (y, clk, wire808, wire807, wire806, wire805);
  output wire [(32'h528):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h10):(1'h0)] wire808;
  input wire signed [(4'hc):(1'h0)] wire807;
  input wire [(3'h4):(1'h0)] wire806;
  input wire signed [(3'h7):(1'h0)] wire805;
  wire signed [(5'h18):(1'h0)] wire851;
  wire signed [(4'hd):(1'h0)] wire850;
  wire [(4'hf):(1'h0)] wire849;
  wire [(5'h11):(1'h0)] wire847;
  wire [(5'h10):(1'h0)] wire846;
  wire signed [(4'h9):(1'h0)] wire845;
  wire signed [(5'h11):(1'h0)] wire839;
  wire [(4'h8):(1'h0)] wire838;
  wire signed [(5'h14):(1'h0)] wire809;
  reg [(5'h14):(1'h0)] reg907 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg903 = (1'h0);
  reg [(5'h11):(1'h0)] reg900 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg899 = (1'h0);
  reg [(4'h8):(1'h0)] reg897 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg895 = (1'h0);
  reg [(5'h15):(1'h0)] reg892 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg891 = (1'h0);
  reg [(4'h9):(1'h0)] reg890 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg889 = (1'h0);
  reg [(4'hb):(1'h0)] reg888 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg887 = (1'h0);
  reg [(5'h16):(1'h0)] reg884 = (1'h0);
  reg [(5'h14):(1'h0)] reg881 = (1'h0);
  reg [(4'ha):(1'h0)] reg877 = (1'h0);
  reg [(3'h7):(1'h0)] reg861 = (1'h0);
  reg [(5'h12):(1'h0)] reg871 = (1'h0);
  reg [(3'h5):(1'h0)] reg870 = (1'h0);
  reg [(4'ha):(1'h0)] reg868 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg865 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg863 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg862 = (1'h0);
  reg [(5'h10):(1'h0)] reg859 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg858 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg857 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg855 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg844 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg843 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg842 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg841 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg837 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg834 = (1'h0);
  reg [(4'h9):(1'h0)] reg833 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg832 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg825 = (1'h0);
  reg [(5'h10):(1'h0)] reg823 = (1'h0);
  reg [(4'hd):(1'h0)] reg822 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg821 = (1'h0);
  reg [(4'hd):(1'h0)] reg820 = (1'h0);
  reg [(4'h9):(1'h0)] reg819 = (1'h0);
  reg [(4'hd):(1'h0)] reg818 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg817 = (1'h0);
  reg [(5'h10):(1'h0)] reg816 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg814 = (1'h0);
  reg [(2'h2):(1'h0)] reg812 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg906 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar905 = (1'h0);
  reg [(4'hd):(1'h0)] reg904 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar902 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg901 = (1'h0);
  reg [(4'hd):(1'h0)] forvar896 = (1'h0);
  reg [(4'ha):(1'h0)] reg898 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg896 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg894 = (1'h0);
  reg [(5'h18):(1'h0)] reg893 = (1'h0);
  reg [(4'ha):(1'h0)] forvar882 = (1'h0);
  reg [(2'h3):(1'h0)] reg886 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg885 = (1'h0);
  reg [(4'he):(1'h0)] reg883 = (1'h0);
  reg [(2'h3):(1'h0)] reg882 = (1'h0);
  reg [(4'h8):(1'h0)] reg880 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg879 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg878 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar876 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar875 = (1'h0);
  reg [(4'h9):(1'h0)] reg874 = (1'h0);
  reg [(5'h16):(1'h0)] reg873 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg872 = (1'h0);
  reg [(4'he):(1'h0)] reg869 = (1'h0);
  reg [(4'h9):(1'h0)] reg867 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg866 = (1'h0);
  reg [(2'h2):(1'h0)] reg864 = (1'h0);
  reg [(2'h3):(1'h0)] forvar861 = (1'h0);
  reg [(3'h5):(1'h0)] reg860 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg856 = (1'h0);
  reg [(5'h12):(1'h0)] forvar854 = (1'h0);
  reg [(5'h12):(1'h0)] reg853 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg852 = (1'h0);
  reg [(2'h2):(1'h0)] reg848 = (1'h0);
  reg [(5'h15):(1'h0)] reg840 = (1'h0);
  reg [(4'hd):(1'h0)] reg815 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar812 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg836 = (1'h0);
  reg [(5'h14):(1'h0)] reg835 = (1'h0);
  reg [(4'h9):(1'h0)] reg831 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg830 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg829 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar828 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg827 = (1'h0);
  reg [(3'h7):(1'h0)] reg826 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg824 = (1'h0);
  reg [(5'h14):(1'h0)] forvar815 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg813 = (1'h0);
  reg signed [(4'he):(1'h0)] reg811 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg810 = (1'h0);
  assign y = {wire851,
                 wire850,
                 wire849,
                 wire847,
                 wire846,
                 wire845,
                 wire839,
                 wire838,
                 wire809,
                 reg907,
                 reg903,
                 reg900,
                 reg899,
                 reg897,
                 reg895,
                 reg892,
                 reg891,
                 reg890,
                 reg889,
                 reg888,
                 reg887,
                 reg884,
                 reg881,
                 reg877,
                 reg861,
                 reg871,
                 reg870,
                 reg868,
                 reg865,
                 reg863,
                 reg862,
                 reg859,
                 reg858,
                 reg857,
                 reg855,
                 reg844,
                 reg843,
                 reg842,
                 reg841,
                 reg837,
                 reg834,
                 reg833,
                 reg832,
                 reg825,
                 reg823,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 reg818,
                 reg817,
                 reg816,
                 reg814,
                 reg812,
                 reg906,
                 forvar905,
                 reg904,
                 forvar902,
                 reg901,
                 forvar896,
                 reg898,
                 reg896,
                 reg894,
                 reg893,
                 forvar882,
                 reg886,
                 reg885,
                 reg883,
                 reg882,
                 reg880,
                 reg879,
                 reg878,
                 forvar876,
                 forvar875,
                 reg874,
                 reg873,
                 reg872,
                 reg869,
                 reg867,
                 reg866,
                 reg864,
                 forvar861,
                 reg860,
                 reg856,
                 forvar854,
                 reg853,
                 reg852,
                 reg848,
                 reg840,
                 reg815,
                 forvar812,
                 reg836,
                 reg835,
                 reg831,
                 reg830,
                 reg829,
                 forvar828,
                 reg827,
                 reg826,
                 reg824,
                 forvar815,
                 reg813,
                 reg811,
                 reg810,
                 (1'h0)};
  assign wire809 = $signed((wire806[(2'h2):(2'h2)] ?
                       (~^$signed($unsigned(wire805))) : $unsigned(wire808[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      if ($signed($unsigned(({(~wire808)} ?
          (&$signed((7'h4a))) : ((wire806 ? (7'h41) : wire808) ?
              $signed(wire807) : $signed(wire807))))))
        begin
          if ((^(wire808 ~^ wire807[(3'h7):(3'h5)])))
            begin
              reg810 = (|wire805[(1'h0):(1'h0)]);
              reg811 = wire806;
            end
          else
            begin
              reg812 <= $signed((~&wire809));
              reg813 = wire808;
              reg814 <= (wire808[(4'hf):(1'h1)] ?
                  reg812[(2'h2):(1'h1)] : (+((wire808[(4'h9):(3'h6)] ?
                      $unsigned(reg813) : wire809) ^ $unsigned({wire805}))));
            end
          for (forvar815 = (1'h0); (forvar815 < (1'h0)); forvar815 = (forvar815 + (1'h1)))
            begin
              reg816 <= (((wire805 ?
                  (8'ha2) : reg813[(1'h1):(1'h0)]) << {reg813[(3'h5):(1'h0)],
                  (~|wire806)}) < $signed(((-{reg810, wire809}) & (|{reg813,
                  wire806}))));
              reg817 <= (~|reg811[(2'h2):(1'h0)]);
              reg818 <= $unsigned(((~(forvar815[(5'h12):(4'hb)] ?
                  (&reg816) : (wire808 ? wire807 : forvar815))) * wire807));
            end
          if ((+reg811[(2'h2):(1'h0)]))
            begin
              reg819 <= wire805;
              reg820 <= wire807;
              reg821 <= reg811[(3'h7):(2'h2)];
              reg822 <= (&reg816);
              reg823 <= wire805;
            end
          else
            begin
              reg824 = {reg813[(3'h5):(3'h4)]};
              reg825 <= (8'ha9);
              reg826 = reg821;
              reg827 = $signed((reg814[(5'h10):(4'h9)] ?
                  $unsigned($signed(((8'haf) ?
                      reg814 : reg822))) : (^~forvar815)));
            end
          for (forvar828 = (1'h0); (forvar828 < (1'h1)); forvar828 = (forvar828 + (1'h1)))
            begin
              reg829 = reg814[(3'h7):(1'h0)];
              reg830 = $signed(reg820[(3'h6):(3'h5)]);
              reg831 = $signed((~^reg811));
              reg832 <= reg830[(2'h3):(2'h3)];
            end
          if ($signed(((((-reg831) ?
              $unsigned((8'hb0)) : reg825[(4'h8):(4'h8)]) > (^~(reg831 ?
              reg824 : reg813))) && ((reg822[(3'h7):(1'h1)] ^ $signed(reg813)) ?
              $unsigned($signed(reg819)) : ((reg814 - (7'h41)) ?
                  (reg826 ? reg814 : (8'hb5)) : (reg832 ? reg811 : (8'ha0)))))))
            begin
              reg833 <= ((reg810 ~^ (wire808 | $unsigned((reg816 ?
                  reg814 : reg819)))) < reg821);
              reg834 <= (~^(~(~&(reg814 & $signed(reg829)))));
              reg835 = reg834[(3'h5):(3'h5)];
              reg836 = (~$signed(wire806));
              reg837 <= ($signed(reg829) > $signed((wire809 ?
                  (^~(reg813 * (8'ha9))) : $signed((^reg822)))));
            end
          else
            begin
              reg835 = $signed((&((reg810[(3'h5):(3'h5)] >>> ((8'ha6) ?
                  (8'ha4) : reg810)) >> (~&(reg837 ? reg820 : (8'hae))))));
              reg836 = ($unsigned(reg824) ?
                  $signed((&$signed(reg814[(4'ha):(3'h7)]))) : reg829[(2'h3):(1'h0)]);
            end
        end
      else
        begin
          reg810 = ((reg822[(4'h9):(3'h7)] ?
                  ((reg819 ?
                      $signed(reg812) : $signed((7'h45))) >= reg823) : reg813[(2'h3):(2'h3)]) ?
              (|$signed({$signed((7'h45))})) : reg835[(4'hf):(3'h7)]);
          reg811 = ($signed(reg821[(4'ha):(3'h7)]) ^~ (reg830[(4'h9):(4'h9)] ?
              $signed($signed($signed(forvar828))) : $signed(reg814[(3'h6):(1'h1)])));
          for (forvar812 = (1'h0); (forvar812 < (1'h0)); forvar812 = (forvar812 + (1'h1)))
            begin
              reg813 = (~^$signed(reg831[(1'h0):(1'h0)]));
              reg815 = $signed((|(reg825[(4'ha):(2'h3)] < (reg834[(3'h7):(1'h0)] >> (wire809 + wire805)))));
              reg824 = (reg827[(1'h0):(1'h0)] == forvar815[(5'h10):(4'h8)]);
              reg826 = $unsigned((&{forvar815}));
            end
        end
    end
  assign wire838 = $unsigned({reg832[(1'h0):(1'h0)],
                       ((~^(wire809 || reg820)) ^~ (&$unsigned(reg820)))});
  assign wire839 = reg823[(3'h6):(3'h6)];
  always
    @(posedge clk) begin
      reg840 = reg812;
    end
  always
    @(posedge clk) begin
      reg841 <= ({$signed(wire839[(1'h1):(1'h0)]),
          $unsigned(reg837[(1'h1):(1'h0)])} << reg832);
      reg842 <= $unsigned((^~((reg822[(1'h1):(1'h1)] ?
              (~&reg817) : $unsigned(wire805)) ?
          (reg834 ~^ reg832) : reg833)));
      reg843 <= (^~$signed($signed((~{wire839, reg818}))));
      reg844 <= (wire807[(4'h9):(3'h5)] ?
          wire808 : (($signed((reg818 ? reg822 : reg834)) ^ (reg818 ?
                  (8'ha4) : (reg832 == reg820))) ?
              wire808[(3'h6):(1'h0)] : (8'h9f)));
    end
  assign wire845 = (reg843 >= $unsigned((-((wire806 ? reg834 : reg821) ?
                       reg841[(5'h11):(4'hb)] : $unsigned(wire807)))));
  assign wire846 = ((wire838 > $signed(($signed(wire805) ?
                           $signed((8'hb9)) : wire809))) ?
                       $signed($unsigned(({reg823} - (reg832 >> reg818)))) : (8'hb1));
  assign wire847 = $unsigned((($signed((reg814 ?
                       wire846 : reg841)) | (!$unsigned(reg817))) > wire809[(2'h3):(1'h0)]));
  always
    @(posedge clk) begin
      reg848 = (!wire806[(3'h4):(1'h1)]);
    end
  assign wire849 = reg821;
  assign wire850 = ({(|wire849[(4'hb):(2'h2)]),
                           $unsigned((wire808[(4'hf):(4'ha)] <= (wire839 ?
                               reg812 : reg812)))} ?
                       (reg837[(2'h2):(1'h1)] << (((|wire807) ?
                           (wire839 >> reg812) : (~|wire809)) ^~ ((wire847 << reg814) ?
                           ((8'ha9) || wire839) : $unsigned(wire805)))) : (($unsigned({wire847}) ?
                           (8'hb4) : $signed(wire849[(2'h3):(2'h3)])) ~^ ($signed((wire807 ?
                           (8'h9f) : reg844)) ^~ reg825)));
  assign wire851 = $unsigned((reg814 - ((((8'h9d) ? wire808 : wire838) ?
                           $unsigned(wire847) : $unsigned(reg844)) ?
                       ({reg820, reg834} ?
                           (~^reg817) : ((8'hba) && reg812)) : $unsigned($signed(wire846)))));
  always
    @(posedge clk) begin
      reg852 = wire808[(4'h9):(1'h1)];
      reg853 = wire847;
      for (forvar854 = (1'h0); (forvar854 < (2'h2)); forvar854 = (forvar854 + (1'h1)))
        begin
          reg855 <= ($unsigned(wire851) ?
              {$unsigned((7'h4a))} : (|($unsigned(reg825[(4'h8):(4'h8)]) ?
                  ($unsigned(reg833) >= reg833) : $signed($signed(wire849)))));
          reg856 = ($unsigned($unsigned(reg833[(2'h3):(2'h2)])) + $signed(wire805));
          reg857 <= (-reg814[(3'h6):(1'h0)]);
          reg858 <= (((($unsigned(wire807) ?
              (wire838 != reg843) : wire845) || ((!wire845) ^ (^wire845))) ^ (^$signed((~&reg833)))) * reg856[(3'h4):(1'h0)]);
          reg859 <= (reg855[(2'h3):(2'h3)] ?
              (|(($signed((8'haf)) >>> {wire807, wire807}) ?
                  (+(wire850 > wire849)) : ({reg855, reg832} ?
                      reg820[(1'h0):(1'h0)] : $unsigned(reg812)))) : $signed(forvar854[(3'h7):(3'h6)]));
        end
      reg860 = (reg859 - reg820);
      if (($signed(reg825[(1'h1):(1'h0)]) ?
          {reg818[(4'hc):(4'hb)], reg822} : $unsigned(reg859)))
        begin
          for (forvar861 = (1'h0); (forvar861 < (2'h2)); forvar861 = (forvar861 + (1'h1)))
            begin
              reg862 <= (reg841 ?
                  reg817 : (wire850 ?
                      ($signed(reg817[(3'h4):(3'h4)]) ?
                          wire806[(1'h1):(1'h1)] : reg820[(3'h4):(3'h4)]) : (~wire807[(2'h2):(2'h2)])));
              reg863 <= $signed({((!(~|reg841)) + $unsigned($unsigned(reg832)))});
            end
          reg864 = $unsigned({(^~$signed(wire809[(4'hb):(4'ha)])),
              reg857[(1'h0):(1'h0)]});
          reg865 <= (-$unsigned($signed($signed((|wire850)))));
          if (({reg814[(2'h2):(1'h0)],
                  (($unsigned(reg819) ?
                      $signed(reg834) : {wire847,
                          reg814}) > $unsigned($unsigned(forvar854)))} ?
              ((((reg823 ? (8'h9c) : reg857) ?
                      (wire809 << (8'ha8)) : (reg823 ? reg865 : reg852)) ?
                  $unsigned({reg837,
                      reg857}) : (~$unsigned((7'h42)))) && wire808[(3'h7):(2'h2)]) : ($unsigned((~&wire806)) ?
                  (~((reg864 ^~ reg860) ^ (reg852 | wire805))) : $signed($unsigned((reg844 ?
                      reg819 : reg843))))))
            begin
              reg866 = wire807;
              reg867 = (^~{$signed(((-forvar861) ~^ (+reg812)))});
              reg868 <= reg833;
            end
          else
            begin
              reg868 <= $signed(forvar854[(3'h7):(3'h6)]);
              reg869 = reg822[(4'hb):(3'h7)];
              reg870 <= (($signed(reg868[(2'h3):(1'h1)]) >= reg822) ?
                  (($signed($signed(reg821)) ^~ $unsigned((^~forvar854))) != ({$signed((7'h4a)),
                      $signed(reg822)} != (reg834 || ((7'h47) > reg823)))) : (reg814[(3'h4):(1'h1)] != (!reg822[(3'h4):(3'h4)])));
              reg871 <= {((((reg843 ? wire809 : reg834) ?
                          (~&reg841) : reg858[(3'h7):(3'h7)]) > $signed($unsigned((8'hb3)))) ?
                      (~&$signed(reg833[(3'h6):(3'h6)])) : reg817),
                  $unsigned((!reg832[(1'h1):(1'h0)]))};
            end
          reg872 = reg812[(2'h2):(1'h1)];
        end
      else
        begin
          reg861 <= (reg870 == {(~wire849), (!$signed(reg812[(1'h1):(1'h1)]))});
          if ($signed(reg820[(3'h5):(2'h3)]))
            begin
              reg864 = (^reg860[(1'h1):(1'h1)]);
              reg866 = (~|(((~(+reg843)) <= $unsigned(reg832)) == $signed(reg855[(3'h4):(2'h2)])));
              reg867 = $unsigned((+((~$unsigned(wire839)) - reg822[(4'h8):(3'h7)])));
            end
          else
            begin
              reg862 <= (7'h43);
              reg864 = $unsigned(reg817[(3'h6):(2'h2)]);
              reg865 <= (|$signed(wire807));
            end
          if ({reg862[(1'h1):(1'h1)]})
            begin
              reg869 = $unsigned($unsigned(((^~reg818) | reg853[(1'h0):(1'h0)])));
              reg870 <= (&($signed(({reg825, reg818} ? wire806 : {wire806})) ?
                  (~&wire849) : ($signed(reg869[(2'h3):(2'h3)]) == $signed($signed(wire806)))));
            end
          else
            begin
              reg868 <= (8'h9f);
            end
        end
    end
  always
    @(posedge clk) begin
      reg873 = $unsigned(($unsigned(($signed(reg832) | reg861[(3'h7):(3'h5)])) ^~ (reg832[(2'h2):(1'h1)] >>> reg834[(4'h9):(1'h0)])));
      reg874 = reg858[(2'h2):(1'h0)];
    end
  always
    @(posedge clk) begin
      for (forvar875 = (1'h0); (forvar875 < (2'h3)); forvar875 = (forvar875 + (1'h1)))
        begin
          for (forvar876 = (1'h0); (forvar876 < (2'h2)); forvar876 = (forvar876 + (1'h1)))
            begin
              reg877 <= reg832[(2'h2):(2'h2)];
              reg878 = (!wire808[(4'h8):(3'h6)]);
              reg879 = $signed({wire847});
              reg880 = ($unsigned($unsigned(($unsigned(wire849) | $unsigned(reg833)))) ~^ {($unsigned(reg832) ?
                      reg879[(2'h3):(1'h1)] : reg843[(1'h1):(1'h0)]),
                  reg870});
            end
        end
      reg881 <= (($signed(wire839[(3'h7):(3'h6)]) & (|(^(+(7'h45))))) ?
          (+(+reg825)) : ((!wire806) ?
              $unsigned((+{(8'hb8)})) : $signed($unsigned(reg865[(5'h10):(1'h0)]))));
      if ({$unsigned({wire845[(3'h7):(3'h4)], (~$signed(reg832))}),
          (-$unsigned(reg837))})
        begin
          if (({reg833,
              ($signed((reg822 ?
                  (8'ha0) : reg868)) >= $signed((reg881 > (8'hb0))))} >= {$signed(reg833),
              (+((reg877 ? reg817 : reg881) <= (~wire849)))}))
            begin
              reg882 = ((!(reg861 << wire850)) >>> ((~(((7'h49) - reg842) ?
                  reg844 : (forvar875 < (8'ha3)))) > $signed((!((8'hac) ?
                  reg841 : reg842)))));
              reg883 = $unsigned(reg870[(2'h3):(1'h0)]);
              reg884 <= (&(~wire847[(3'h7):(2'h2)]));
              reg885 = reg832;
              reg886 = (-{({(&reg885)} >>> reg868[(3'h5):(1'h0)])});
            end
          else
            begin
              reg882 = (~(reg832 ?
                  (~((+reg865) ?
                      (~&reg879) : $unsigned(reg868))) : (reg843[(3'h4):(3'h4)] ?
                      $unsigned((reg818 >> reg841)) : $unsigned((reg858 ?
                          reg822 : wire805)))));
              reg884 <= {reg883[(3'h5):(1'h0)]};
              reg885 = reg882;
            end
          reg887 <= {$signed($unsigned(reg857)), wire809[(4'hf):(3'h5)]};
          reg888 <= (~|$signed((reg825 ^ ((^~reg882) ?
              reg884 : ((8'h9c) ? reg812 : reg879)))));
        end
      else
        begin
          for (forvar882 = (1'h0); (forvar882 < (3'h4)); forvar882 = (forvar882 + (1'h1)))
            begin
              reg884 <= $unsigned($signed(reg818));
              reg887 <= ($signed(reg812) ?
                  reg859[(4'he):(4'h8)] : $signed(reg843[(3'h4):(1'h0)]));
              reg888 <= ($unsigned((!((+reg883) ?
                      reg832[(2'h2):(1'h0)] : reg841[(3'h7):(1'h1)]))) ?
                  $signed(($signed((reg832 ^ reg825)) && ((reg861 ^~ reg878) ?
                      wire809[(4'ha):(1'h0)] : (wire808 ?
                          (7'h44) : reg886)))) : $unsigned((8'hbc)));
            end
          reg889 <= (+reg888[(1'h0):(1'h0)]);
          reg890 <= (($unsigned(($unsigned((8'hb5)) ?
              (reg859 ?
                  reg884 : wire805) : {reg844})) != $unsigned($signed($signed(reg888)))) * $signed($unsigned($signed((forvar875 ?
              reg871 : reg865)))));
          reg891 <= wire847[(2'h2):(2'h2)];
          reg892 <= $signed(({(reg880[(1'h1):(1'h1)] ?
                  reg822[(3'h6):(3'h6)] : {reg877, (7'h40)}),
              ($unsigned(forvar882) ?
                  $unsigned(reg817) : $signed(reg881))} && (reg882[(2'h3):(1'h0)] ?
              $signed((|reg863)) : ((^(8'hb0)) ?
                  (~|(8'ha1)) : reg819[(2'h3):(1'h1)]))));
        end
      reg893 = $signed(reg884);
      if ((!{$signed((7'h48))}))
        begin
          reg894 = ((8'h9f) == reg885);
          if ((&((reg817 ?
              $unsigned(reg823) : ({wire851, reg861} ?
                  reg889 : reg819[(2'h2):(2'h2)])) ^ reg832[(2'h2):(1'h1)])))
            begin
              reg895 <= reg812;
              reg896 = (^{reg814[(1'h1):(1'h1)],
                  ($signed((reg865 ? reg865 : reg833)) * {$signed(reg837),
                      $signed(reg890)})});
              reg897 <= (reg862 <= reg821);
              reg898 = {reg887,
                  $unsigned((((8'hb0) <<< {reg814, reg859}) ?
                      $unsigned($signed(reg894)) : reg817[(3'h4):(3'h4)]))};
            end
          else
            begin
              reg896 = forvar876[(4'hd):(4'h9)];
            end
          if (($unsigned(reg883[(4'hd):(3'h6)]) && $signed($signed($unsigned({reg886,
              (8'haa)})))))
            begin
              reg899 <= $unsigned(({$signed({(8'hb3)})} ^~ $unsigned(forvar875[(3'h5):(2'h3)])));
            end
          else
            begin
              reg899 <= $signed((^(~&$unsigned(reg841))));
            end
          reg900 <= reg899[(4'hd):(3'h6)];
        end
      else
        begin
          reg895 <= $unsigned(reg888);
          for (forvar896 = (1'h0); (forvar896 < (3'h4)); forvar896 = (forvar896 + (1'h1)))
            begin
              reg897 <= forvar896[(1'h1):(1'h0)];
              reg899 <= {(-((~&(reg833 ? reg890 : (8'hb2))) ?
                      reg865 : ((wire845 * reg881) ?
                          wire846[(3'h5):(3'h4)] : $unsigned(reg833))))};
              reg901 = (reg834[(4'ha):(2'h3)] || $signed(((~^((8'ha1) | reg894)) ?
                  (^~reg822[(4'hc):(4'h8)]) : $signed((reg834 == reg897)))));
            end
          for (forvar902 = (1'h0); (forvar902 < (2'h3)); forvar902 = (forvar902 + (1'h1)))
            begin
              reg903 <= (reg822 ?
                  $signed((reg844 ?
                      $signed(reg892) : reg862)) : reg888[(4'h8):(3'h5)]);
            end
          reg904 = reg903[(3'h7):(1'h0)];
          for (forvar905 = (1'h0); (forvar905 < (2'h3)); forvar905 = (forvar905 + (1'h1)))
            begin
              reg906 = $signed($unsigned((~forvar905)));
              reg907 <= $signed((^~reg823[(4'ha):(3'h6)]));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module578
#(parameter param737 = ((((!((8'ha1) ? (8'hb5) : (8'ha5))) ? (((8'ha6) ? (8'ha9) : (8'hbe)) ? ((7'h40) ? (8'h9e) : (8'h9c)) : (^~(7'h41))) : (((8'hb7) ? (8'h9c) : (8'ha9)) <= (|(8'ha8)))) ? ((((8'ha4) ? (8'ha0) : (7'h42)) ? ((8'hbe) ? (8'ha5) : (7'h42)) : ((7'h40) ? (8'hb9) : (8'h9f))) ? ((~&(8'hb0)) ? ((8'hae) <<< (8'hab)) : (8'ha1)) : (((7'h49) & (8'hb3)) ? ((8'hb6) ? (8'ha5) : (8'hb7)) : ((8'h9d) ? (8'h9d) : (7'h45)))) : (((^(8'hbf)) ~^ {(8'haf)}) ? (~|(^~(7'h44))) : (((7'h46) & (8'ha0)) * (~(8'hab))))) ? ({((^~(7'h44)) ? ((8'hb7) ^ (8'hb7)) : (~&(8'ha2))), (((8'ha6) > (8'hac)) ? ((8'ha5) == (8'ha5)) : (~(8'hb3)))} + {((~(7'h44)) <= {(8'ha7)})}) : (+(^{((8'hac) + (7'h49)), (^(8'hb2))}))))
(y, clk, wire583, wire582, wire581, wire580, wire579);
  output wire [(32'h856):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire583;
  input wire signed [(5'h13):(1'h0)] wire582;
  input wire signed [(4'h8):(1'h0)] wire581;
  input wire signed [(4'ha):(1'h0)] wire580;
  input wire signed [(5'h12):(1'h0)] wire579;
  wire signed [(4'he):(1'h0)] wire736;
  wire [(4'hb):(1'h0)] wire735;
  wire signed [(4'hf):(1'h0)] wire734;
  wire signed [(4'hb):(1'h0)] wire702;
  wire [(5'h18):(1'h0)] wire701;
  wire [(5'h17):(1'h0)] wire700;
  wire [(5'h10):(1'h0)] wire648;
  wire signed [(5'h14):(1'h0)] wire647;
  wire signed [(2'h3):(1'h0)] wire618;
  wire [(3'h5):(1'h0)] wire617;
  wire signed [(5'h11):(1'h0)] wire591;
  wire [(3'h6):(1'h0)] wire585;
  wire [(4'h8):(1'h0)] wire584;
  reg signed [(5'h18):(1'h0)] reg733 = (1'h0);
  reg [(3'h6):(1'h0)] reg732 = (1'h0);
  reg [(5'h14):(1'h0)] reg729 = (1'h0);
  reg [(5'h16):(1'h0)] reg725 = (1'h0);
  reg [(5'h11):(1'h0)] reg724 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg723 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg717 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg716 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg715 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg711 = (1'h0);
  reg [(4'he):(1'h0)] reg710 = (1'h0);
  reg [(3'h7):(1'h0)] reg708 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg699 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg698 = (1'h0);
  reg [(4'he):(1'h0)] reg697 = (1'h0);
  reg [(3'h5):(1'h0)] reg683 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg689 = (1'h0);
  reg [(5'h14):(1'h0)] reg686 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg684 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg682 = (1'h0);
  reg [(3'h5):(1'h0)] reg675 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg674 = (1'h0);
  reg [(4'hb):(1'h0)] reg671 = (1'h0);
  reg [(4'h8):(1'h0)] reg670 = (1'h0);
  reg [(5'h17):(1'h0)] reg669 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg668 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg664 = (1'h0);
  reg [(3'h6):(1'h0)] reg660 = (1'h0);
  reg [(5'h17):(1'h0)] reg659 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg655 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg654 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg649 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg646 = (1'h0);
  reg [(3'h4):(1'h0)] reg645 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg642 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg641 = (1'h0);
  reg signed [(4'he):(1'h0)] reg640 = (1'h0);
  reg [(2'h3):(1'h0)] reg637 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg634 = (1'h0);
  reg signed [(4'he):(1'h0)] reg632 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg631 = (1'h0);
  reg [(5'h13):(1'h0)] reg630 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg629 = (1'h0);
  reg signed [(4'he):(1'h0)] reg626 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg623 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg616 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg614 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg613 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg612 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg609 = (1'h0);
  reg [(5'h11):(1'h0)] reg607 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg602 = (1'h0);
  reg [(4'hb):(1'h0)] reg596 = (1'h0);
  reg [(4'h8):(1'h0)] reg594 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg593 = (1'h0);
  reg [(5'h18):(1'h0)] reg590 = (1'h0);
  reg [(5'h16):(1'h0)] reg586 = (1'h0);
  reg [(3'h4):(1'h0)] reg731 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg730 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg728 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg727 = (1'h0);
  reg [(4'hf):(1'h0)] reg726 = (1'h0);
  reg [(5'h10):(1'h0)] reg722 = (1'h0);
  reg [(5'h14):(1'h0)] reg721 = (1'h0);
  reg [(5'h11):(1'h0)] reg720 = (1'h0);
  reg [(4'hb):(1'h0)] reg719 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar718 = (1'h0);
  reg [(5'h14):(1'h0)] reg714 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg713 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar712 = (1'h0);
  reg [(4'ha):(1'h0)] reg709 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg707 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg706 = (1'h0);
  reg [(2'h3):(1'h0)] reg705 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg704 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar703 = (1'h0);
  reg [(4'ha):(1'h0)] reg696 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg695 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar694 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg693 = (1'h0);
  reg [(4'h8):(1'h0)] reg692 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar691 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar686 = (1'h0);
  reg [(3'h4):(1'h0)] reg685 = (1'h0);
  reg [(3'h6):(1'h0)] forvar675 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg673 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg690 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg688 = (1'h0);
  reg [(3'h4):(1'h0)] reg687 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar685 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar683 = (1'h0);
  reg [(5'h12):(1'h0)] reg681 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg680 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg679 = (1'h0);
  reg [(3'h7):(1'h0)] reg678 = (1'h0);
  reg signed [(4'he):(1'h0)] reg677 = (1'h0);
  reg [(4'hd):(1'h0)] reg676 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar673 = (1'h0);
  reg [(3'h6):(1'h0)] reg672 = (1'h0);
  reg [(5'h10):(1'h0)] forvar667 = (1'h0);
  reg [(4'hf):(1'h0)] forvar666 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg665 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg663 = (1'h0);
  reg [(5'h17):(1'h0)] reg662 = (1'h0);
  reg [(5'h13):(1'h0)] reg661 = (1'h0);
  reg [(5'h12):(1'h0)] reg658 = (1'h0);
  reg [(5'h17):(1'h0)] forvar657 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg656 = (1'h0);
  reg [(4'he):(1'h0)] reg653 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg652 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg651 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar650 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg644 = (1'h0);
  reg [(4'hb):(1'h0)] reg643 = (1'h0);
  reg signed [(4'he):(1'h0)] reg639 = (1'h0);
  reg [(5'h18):(1'h0)] forvar638 = (1'h0);
  reg [(4'hb):(1'h0)] reg636 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg635 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg633 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar628 = (1'h0);
  reg [(5'h17):(1'h0)] forvar627 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg625 = (1'h0);
  reg [(3'h6):(1'h0)] reg624 = (1'h0);
  reg [(4'hd):(1'h0)] reg622 = (1'h0);
  reg [(5'h15):(1'h0)] reg621 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar620 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg619 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg615 = (1'h0);
  reg [(5'h16):(1'h0)] forvar601 = (1'h0);
  reg [(3'h5):(1'h0)] forvar611 = (1'h0);
  reg [(4'he):(1'h0)] reg610 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg608 = (1'h0);
  reg [(4'hb):(1'h0)] forvar606 = (1'h0);
  reg [(5'h11):(1'h0)] reg605 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg604 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg603 = (1'h0);
  reg signed [(4'he):(1'h0)] reg601 = (1'h0);
  reg [(5'h15):(1'h0)] reg600 = (1'h0);
  reg [(2'h3):(1'h0)] reg599 = (1'h0);
  reg [(4'h9):(1'h0)] reg598 = (1'h0);
  reg signed [(4'he):(1'h0)] reg597 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg595 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar592 = (1'h0);
  reg [(4'h8):(1'h0)] reg589 = (1'h0);
  reg signed [(4'he):(1'h0)] reg588 = (1'h0);
  reg [(4'hc):(1'h0)] forvar587 = (1'h0);
  assign y = {wire736,
                 wire735,
                 wire734,
                 wire702,
                 wire701,
                 wire700,
                 wire648,
                 wire647,
                 wire618,
                 wire617,
                 wire591,
                 wire585,
                 wire584,
                 reg733,
                 reg732,
                 reg729,
                 reg725,
                 reg724,
                 reg723,
                 reg717,
                 reg716,
                 reg715,
                 reg711,
                 reg710,
                 reg708,
                 reg699,
                 reg698,
                 reg697,
                 reg683,
                 reg689,
                 reg686,
                 reg684,
                 reg682,
                 reg675,
                 reg674,
                 reg671,
                 reg670,
                 reg669,
                 reg668,
                 reg664,
                 reg660,
                 reg659,
                 reg655,
                 reg654,
                 reg649,
                 reg646,
                 reg645,
                 reg642,
                 reg641,
                 reg640,
                 reg637,
                 reg634,
                 reg632,
                 reg631,
                 reg630,
                 reg629,
                 reg626,
                 reg623,
                 reg616,
                 reg614,
                 reg613,
                 reg612,
                 reg609,
                 reg607,
                 reg602,
                 reg596,
                 reg594,
                 reg593,
                 reg590,
                 reg586,
                 reg731,
                 reg730,
                 reg728,
                 reg727,
                 reg726,
                 reg722,
                 reg721,
                 reg720,
                 reg719,
                 forvar718,
                 reg714,
                 reg713,
                 forvar712,
                 reg709,
                 reg707,
                 reg706,
                 reg705,
                 reg704,
                 forvar703,
                 reg696,
                 reg695,
                 forvar694,
                 reg693,
                 reg692,
                 forvar691,
                 forvar686,
                 reg685,
                 forvar675,
                 reg673,
                 reg690,
                 reg688,
                 reg687,
                 forvar685,
                 forvar683,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 reg677,
                 reg676,
                 forvar673,
                 reg672,
                 forvar667,
                 forvar666,
                 reg665,
                 reg663,
                 reg662,
                 reg661,
                 reg658,
                 forvar657,
                 reg656,
                 reg653,
                 reg652,
                 reg651,
                 forvar650,
                 reg644,
                 reg643,
                 reg639,
                 forvar638,
                 reg636,
                 reg635,
                 reg633,
                 forvar628,
                 forvar627,
                 reg625,
                 reg624,
                 reg622,
                 reg621,
                 forvar620,
                 reg619,
                 reg615,
                 forvar601,
                 forvar611,
                 reg610,
                 reg608,
                 forvar606,
                 reg605,
                 reg604,
                 reg603,
                 reg601,
                 reg600,
                 reg599,
                 reg598,
                 reg597,
                 reg595,
                 forvar592,
                 reg589,
                 reg588,
                 forvar587,
                 (1'h0)};
  assign wire584 = ((-wire580[(4'ha):(3'h5)]) ~^ wire580);
  assign wire585 = wire580[(3'h5):(1'h1)];
  always
    @(posedge clk) begin
      reg586 <= (~^(|(8'h9d)));
      for (forvar587 = (1'h0); (forvar587 < (2'h3)); forvar587 = (forvar587 + (1'h1)))
        begin
          reg588 = ($unsigned($unsigned((~&reg586))) && wire579[(3'h4):(1'h1)]);
          reg589 = reg586[(1'h0):(1'h0)];
        end
      reg590 <= $signed(wire585);
    end
  assign wire591 = $signed(wire581[(4'h8):(1'h0)]);
  always
    @(posedge clk) begin
      for (forvar592 = (1'h0); (forvar592 < (2'h2)); forvar592 = (forvar592 + (1'h1)))
        begin
          if (reg590)
            begin
              reg593 <= wire581;
              reg594 <= $unsigned(((-$signed((reg590 ?
                  wire585 : reg590))) >>> $signed(reg586)));
            end
          else
            begin
              reg595 = $signed({$unsigned({(reg590 - wire585), forvar592}),
                  reg586[(3'h6):(3'h5)]});
              reg596 <= ($unsigned(((7'h45) ?
                  (|wire580) : reg594)) << $unsigned({reg593,
                  $signed(wire581[(2'h3):(2'h3)])}));
              reg597 = reg594;
              reg598 = wire582;
              reg599 = (forvar592 ?
                  ($unsigned(wire579) || $signed((reg597 ?
                      reg586 : $signed(wire583)))) : (+wire584));
            end
          reg600 = $signed($signed(reg599[(1'h1):(1'h1)]));
        end
      if ($signed((~^$signed({$unsigned(wire585)}))))
        begin
          if (reg594[(2'h2):(1'h1)])
            begin
              reg601 = reg597;
              reg602 <= (reg597 ?
                  reg593[(1'h1):(1'h0)] : wire583[(1'h0):(1'h0)]);
            end
          else
            begin
              reg601 = reg600;
              reg603 = $unsigned(reg590);
            end
          reg604 = ($unsigned((($signed(reg598) ?
                  {wire585} : $signed(wire581)) ?
              (reg590 <= (reg599 ?
                  wire585 : reg590)) : wire580)) + $signed((|(reg603[(2'h2):(1'h1)] >>> $unsigned((7'h44))))));
          reg605 = wire579;
          for (forvar606 = (1'h0); (forvar606 < (2'h2)); forvar606 = (forvar606 + (1'h1)))
            begin
              reg607 <= $signed(forvar606);
              reg608 = (~$unsigned(($unsigned((reg599 >= (8'hb5))) ^~ wire582[(2'h2):(1'h0)])));
              reg609 <= $signed($signed(((!(reg596 + reg590)) ?
                  (+(!wire584)) : forvar592)));
              reg610 = ((8'ha9) ?
                  reg609 : ($unsigned($signed($unsigned((8'hbf)))) != reg598[(4'h8):(3'h6)]));
            end
          for (forvar611 = (1'h0); (forvar611 < (2'h3)); forvar611 = (forvar611 + (1'h1)))
            begin
              reg612 <= (reg594[(2'h2):(1'h1)] >>> wire582);
              reg613 <= wire580;
            end
        end
      else
        begin
          for (forvar601 = (1'h0); (forvar601 < (1'h0)); forvar601 = (forvar601 + (1'h1)))
            begin
              reg602 <= reg597;
            end
          reg603 = ($unsigned(reg586[(4'ha):(3'h6)]) ?
              (^(($unsigned(reg607) && $signed(wire591)) ^ reg602)) : wire591);
        end
      reg614 <= (reg604[(4'hb):(3'h7)] ?
          (($unsigned((-(7'h4a))) > $signed((forvar592 ?
              reg601 : forvar606))) && ($signed((7'h43)) >>> (!$signed(forvar592)))) : $unsigned((&$unsigned($signed((8'hb3))))));
      reg615 = $unsigned((|$signed((((8'ha9) == reg586) ?
          (~|forvar611) : (wire584 ? (8'haf) : wire581)))));
    end
  always
    @(posedge clk) begin
      reg616 <= $signed(reg590[(1'h1):(1'h1)]);
    end
  assign wire617 = $signed($signed(reg586[(4'ha):(4'h9)]));
  assign wire618 = $signed($unsigned($unsigned($unsigned(reg614))));
  always
    @(posedge clk) begin
      reg619 = reg602[(4'he):(4'hc)];
      for (forvar620 = (1'h0); (forvar620 < (2'h2)); forvar620 = (forvar620 + (1'h1)))
        begin
          if ((~$unsigned((($unsigned(reg596) ?
                  (wire579 ? reg594 : (8'hac)) : $signed(wire585)) ?
              $unsigned((+reg614)) : $unsigned((reg593 ? reg609 : reg590))))))
            begin
              reg621 = ((|($unsigned(reg607[(3'h4):(2'h2)]) ?
                  wire581[(1'h0):(1'h0)] : reg590)) < $signed(reg614));
              reg622 = (((&((reg609 >= forvar620) ?
                          $signed(reg586) : forvar620)) ?
                      (reg594[(1'h1):(1'h1)] ~^ (~|((7'h49) ?
                          wire584 : wire582))) : ((wire580 ?
                          ((7'h40) != reg613) : (reg593 ?
                              reg614 : (7'h43))) <= (~^{forvar620}))) ?
                  ($unsigned((~|(wire581 * reg590))) ?
                      (^~$signed($unsigned(wire582))) : (8'ha1)) : (($signed(wire583) != (~|(~(8'hb6)))) ~^ $signed(((wire583 * (7'h49)) == $unsigned(wire585)))));
            end
          else
            begin
              reg621 = ($signed((!reg613[(3'h7):(1'h0)])) + reg593);
            end
          reg623 <= wire583[(3'h4):(2'h2)];
          reg624 = ($signed($unsigned($unsigned((reg619 && wire582)))) ?
              $unsigned($unsigned($unsigned($signed((8'ha4))))) : (reg586[(1'h1):(1'h0)] ?
                  $signed($signed($unsigned(wire582))) : $signed(wire617[(2'h3):(2'h2)])));
          if ($signed((^~wire579)))
            begin
              reg625 = reg594;
              reg626 <= $unsigned((wire581 <= wire579[(3'h6):(3'h4)]));
            end
          else
            begin
              reg625 = $signed(($signed((^~forvar620)) != (((~&reg621) << $signed(wire617)) << ((wire582 ^~ reg624) ^ reg612[(5'h16):(3'h4)]))));
            end
        end
      for (forvar627 = (1'h0); (forvar627 < (3'h4)); forvar627 = (forvar627 + (1'h1)))
        begin
          for (forvar628 = (1'h0); (forvar628 < (1'h1)); forvar628 = (forvar628 + (1'h1)))
            begin
              reg629 <= (~$signed((&(|$unsigned(forvar627)))));
              reg630 <= reg616[(1'h0):(1'h0)];
              reg631 <= (|(({(reg619 ? reg602 : reg623)} << ((wire617 ?
                      wire584 : wire591) < wire617)) ?
                  ((|(^~reg619)) ^ reg586[(4'ha):(3'h4)]) : (~|$signed((~reg622)))));
              reg632 <= ({((~^{reg621}) || $unsigned((+wire579)))} ?
                  $unsigned(reg625[(1'h1):(1'h1)]) : ($signed(((reg607 ^ (8'ha6)) ?
                      reg593 : (forvar628 <= reg609))) & (~|({reg623, wire583} ?
                      $signed(forvar620) : (reg594 ? reg607 : reg586)))));
              reg633 = wire618[(1'h1):(1'h0)];
            end
          if ({reg619[(2'h3):(1'h1)],
              $signed((wire618 ? $signed({(8'hbf), reg594}) : reg631))})
            begin
              reg634 <= (^~(reg614 ? {reg586} : reg625[(2'h2):(2'h2)]));
            end
          else
            begin
              reg635 = (wire591 && reg624);
              reg636 = (|(8'had));
              reg637 <= reg633;
            end
          for (forvar638 = (1'h0); (forvar638 < (2'h2)); forvar638 = (forvar638 + (1'h1)))
            begin
              reg639 = $signed(reg625);
            end
          reg640 <= (+$unsigned((~^(|(forvar627 >>> wire591)))));
          if ($signed({reg634}))
            begin
              reg641 <= reg624;
              reg642 <= (8'hb8);
            end
          else
            begin
              reg643 = $signed({reg614[(1'h1):(1'h1)],
                  (|$unsigned({reg640, wire591}))});
              reg644 = (~^reg636[(4'h8):(4'h8)]);
              reg645 <= (reg593[(3'h6):(1'h1)] != ((8'hb9) ?
                  $signed({(reg642 != (8'hab))}) : (~^(~^(forvar638 ?
                      wire618 : wire584)))));
              reg646 <= (~&((~&(reg636[(1'h0):(1'h0)] ?
                  {(8'had), reg642} : ((8'hbe) ?
                      reg619 : reg622))) >>> $unsigned(forvar620)));
            end
        end
    end
  assign wire647 = (reg602 >> (7'h49));
  assign wire648 = (reg594 ?
                       ({$unsigned(((7'h47) >> reg637))} ?
                           {(reg645[(1'h0):(1'h0)] ?
                                   $unsigned(reg594) : $unsigned((8'hb7))),
                               wire582[(5'h13):(4'hc)]} : (-reg641[(5'h10):(1'h0)])) : (($signed((&reg586)) ?
                           {(8'hbd),
                               reg634[(5'h14):(4'hb)]} : $signed((reg586 ^ (7'h44)))) && wire581));
  always
    @(posedge clk) begin
      reg649 <= (~$unsigned(reg623));
    end
  always
    @(posedge clk) begin
      for (forvar650 = (1'h0); (forvar650 < (3'h4)); forvar650 = (forvar650 + (1'h1)))
        begin
          reg651 = wire647[(3'h4):(2'h3)];
          reg652 = $unsigned(wire579[(5'h12):(5'h12)]);
          reg653 = reg632[(3'h4):(1'h1)];
          reg654 <= wire581;
        end
      reg655 <= ($unsigned((|$unsigned(wire617))) < $unsigned({($unsigned(wire647) ?
              (reg609 ^~ reg613) : (wire580 ? wire648 : (8'ha4)))}));
      reg656 = (^({$signed({reg655}), (|reg623)} < reg653[(4'hb):(4'h8)]));
      for (forvar657 = (1'h0); (forvar657 < (1'h0)); forvar657 = (forvar657 + (1'h1)))
        begin
          reg658 = (-$signed(({{reg607, reg607}, (reg654 ? (8'hbf) : (8'ha4))} ?
              $signed((reg609 ? reg613 : (8'hbf))) : $unsigned((~^reg634)))));
          if ($unsigned(wire581))
            begin
              reg659 <= (~wire591[(2'h2):(2'h2)]);
              reg660 <= reg655[(5'h10):(4'hd)];
            end
          else
            begin
              reg661 = reg602;
              reg662 = reg632[(4'hd):(3'h5)];
              reg663 = (^~($unsigned({(^~reg642),
                      (forvar650 ? reg616 : reg593)}) ?
                  $unsigned(reg662) : ((reg631 ^~ (^~reg594)) >>> reg661)));
              reg664 <= (+({$signed((8'hbc))} && ($unsigned(reg637) ?
                  $unsigned((reg629 * reg616)) : wire583[(1'h0):(1'h0)])));
              reg665 = (((7'h4a) - reg640) ?
                  {{((7'h48) <= $signed(reg614)), $signed({(8'hb5), reg640})},
                      ($signed($signed(reg623)) ?
                          reg614 : {(wire585 <<< reg616)})} : $unsigned(reg653));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar666 = (1'h0); (forvar666 < (1'h1)); forvar666 = (forvar666 + (1'h1)))
        begin
          for (forvar667 = (1'h0); (forvar667 < (1'h0)); forvar667 = (forvar667 + (1'h1)))
            begin
              reg668 <= reg607;
              reg669 <= $unsigned($unsigned((reg629[(2'h3):(2'h3)] ^ reg630[(4'h8):(1'h1)])));
            end
          reg670 <= (~|(8'h9e));
          reg671 <= $unsigned($signed(wire647[(4'hf):(4'h8)]));
        end
      reg672 = ((7'h4a) >= (((-reg607) - ($unsigned(reg626) ?
              {reg614} : reg649)) ?
          $unsigned(($unsigned(reg614) ?
              {reg614} : (8'hb7))) : wire591[(3'h6):(3'h5)]));
      if ({wire581[(3'h5):(1'h0)],
          (forvar666 == ($signed({reg632}) >> (reg593 >= $signed(reg631))))})
        begin
          for (forvar673 = (1'h0); (forvar673 < (2'h3)); forvar673 = (forvar673 + (1'h1)))
            begin
              reg674 <= (~|$unsigned(((reg616[(3'h7):(2'h3)] ?
                      $signed((8'hbf)) : wire591[(1'h0):(1'h0)]) ?
                  ($unsigned((8'hbc)) ?
                      $signed(reg642) : reg672[(3'h6):(3'h6)]) : $signed(reg641[(4'h8):(3'h7)]))));
              reg675 <= $signed(wire585);
              reg676 = (forvar666 != {{$unsigned((reg623 ? wire618 : (8'ha9))),
                      (^{reg590, forvar673})}});
              reg677 = reg637;
            end
          if (((($unsigned((reg642 ? wire585 : reg645)) ?
                  $unsigned(reg607) : reg607) ?
              reg634[(2'h3):(2'h2)] : $unsigned({((8'hb5) >= reg640),
                  {reg649}})) < ((~^(~&$signed(wire583))) ?
              $signed((reg593[(4'he):(4'hc)] > (~^reg634))) : reg664)))
            begin
              reg678 = {(~($unsigned((-reg640)) ?
                      reg642[(3'h4):(2'h2)] : (-(~|reg613)))),
                  (7'h48)};
              reg679 = $signed(reg674[(3'h6):(3'h5)]);
              reg680 = (((($signed(wire583) ^~ reg642) >= $unsigned($signed(reg637))) ?
                      ($unsigned(wire618[(2'h3):(1'h1)]) == ($signed(forvar666) ?
                          $unsigned(reg645) : $signed((8'hb4)))) : ((~^(forvar667 ?
                              (7'h47) : reg614)) ?
                          wire584[(3'h5):(1'h1)] : ($signed(wire618) | $signed(reg674)))) ?
                  (8'h9f) : $unsigned(((-(reg676 ?
                      (8'ha1) : forvar666)) & wire647[(3'h6):(2'h3)])));
              reg681 = ($unsigned(($unsigned((wire618 - reg672)) ?
                      ({reg630} * reg586[(3'h6):(3'h6)]) : $signed((~(8'hb8))))) ?
                  $unsigned((reg637 | $signed((reg672 ?
                      reg613 : reg645)))) : reg669);
            end
          else
            begin
              reg682 <= (^((8'hbe) > reg641[(3'h7):(3'h4)]));
            end
          for (forvar683 = (1'h0); (forvar683 < (3'h4)); forvar683 = (forvar683 + (1'h1)))
            begin
              reg684 <= ({$unsigned((^{(8'hb2)})),
                  (reg668[(3'h5):(1'h1)] ?
                      $unsigned(wire591[(4'hc):(4'h9)]) : forvar666)} > reg670);
            end
          for (forvar685 = (1'h0); (forvar685 < (2'h3)); forvar685 = (forvar685 + (1'h1)))
            begin
              reg686 <= $signed(wire583[(1'h1):(1'h1)]);
              reg687 = reg645;
              reg688 = reg675[(1'h0):(1'h0)];
              reg689 <= wire584;
            end
          reg690 = (~^(((~^reg586) != $signed(((7'h44) ?
              reg602 : forvar666))) < (~^($unsigned(reg596) ?
              (8'ha9) : (reg682 ? (8'hbe) : reg614)))));
        end
      else
        begin
          reg673 = reg686[(4'hd):(2'h3)];
          reg674 <= {reg596};
          for (forvar675 = (1'h0); (forvar675 < (1'h1)); forvar675 = (forvar675 + (1'h1)))
            begin
              reg682 <= $unsigned((^~reg642));
              reg683 <= {(((^~reg594) ?
                          ((reg645 ?
                              reg616 : (8'h9f)) ^~ (-reg670)) : wire581) ?
                      $signed(reg689) : ($signed($signed(reg637)) ^ ((~|reg590) * (~^(8'h9e))))),
                  ($signed($signed(forvar673[(4'hb):(3'h4)])) >= {forvar673})};
              reg684 <= reg645;
              reg685 = ((8'ha9) ?
                  ((reg649[(3'h5):(1'h1)] & (~reg672[(1'h0):(1'h0)])) - $signed(((reg613 ?
                      reg671 : forvar685) * $unsigned(wire591)))) : $signed(($signed((reg640 ?
                      forvar667 : reg632)) ^~ (wire579 > $signed(reg634)))));
            end
          for (forvar686 = (1'h0); (forvar686 < (2'h3)); forvar686 = (forvar686 + (1'h1)))
            begin
              reg687 = reg649;
            end
        end
      for (forvar691 = (1'h0); (forvar691 < (1'h1)); forvar691 = (forvar691 + (1'h1)))
        begin
          reg692 = $unsigned(({(wire579[(3'h5):(3'h4)] && $signed(wire579)),
              $unsigned((-reg590))} >= $unsigned((|wire618))));
          reg693 = {$signed(({(+reg672), (~^reg676)} <= reg670[(3'h5):(1'h1)])),
              (~^reg678)};
          for (forvar694 = (1'h0); (forvar694 < (2'h2)); forvar694 = (forvar694 + (1'h1)))
            begin
              reg695 = (wire582 ?
                  $unsigned({wire585, wire582}) : $signed((((reg655 ?
                              reg607 : wire591) ?
                          $unsigned((8'hb9)) : (forvar694 && (8'hbc))) ?
                      (reg642[(3'h7):(1'h0)] * reg634[(5'h15):(5'h12)]) : ($unsigned((7'h41)) ?
                          $signed((8'ha7)) : reg634[(4'hd):(2'h2)]))));
              reg696 = ($unsigned(($unsigned(wire647) && wire585[(2'h3):(2'h2)])) ?
                  reg654 : $unsigned((reg673[(3'h5):(3'h4)] >= {(8'ha8)})));
              reg697 <= (reg655 ?
                  reg692[(1'h0):(1'h0)] : {$signed(reg596),
                      ($signed(forvar685) ?
                          reg626 : forvar691[(1'h0):(1'h0)])});
              reg698 <= reg690[(5'h10):(4'hd)];
            end
          reg699 <= (wire591[(1'h0):(1'h0)] * (reg664[(4'h8):(3'h6)] ?
              (~|$unsigned($signed((8'h9e)))) : reg641));
        end
    end
  assign wire700 = (^((wire581[(2'h2):(2'h2)] ^~ $unsigned({(8'ha9)})) > reg697));
  assign wire701 = reg590[(4'h8):(1'h0)];
  assign wire702 = $unsigned((reg699[(5'h11):(4'hd)] > (~&reg609)));
  always
    @(posedge clk) begin
      for (forvar703 = (1'h0); (forvar703 < (2'h2)); forvar703 = (forvar703 + (1'h1)))
        begin
          reg704 = ((^reg671[(4'ha):(4'ha)]) ?
              (&((^$signed(reg590)) ?
                  reg645 : ($signed((7'h45)) ?
                      reg697[(2'h2):(1'h0)] : $unsigned(reg640)))) : (^~($signed(reg671[(1'h0):(1'h0)]) << $signed((reg614 >= (8'hbd))))));
          if ($signed((wire584 < $signed($unsigned(reg616)))))
            begin
              reg705 = (^(!(&reg594[(3'h4):(2'h2)])));
              reg706 = reg629[(1'h0):(1'h0)];
              reg707 = ((reg660 ?
                      $signed($unsigned(reg683[(3'h5):(1'h1)])) : $unsigned(($signed((7'h40)) - reg607))) ?
                  $signed(wire702) : reg669[(5'h13):(2'h3)]);
              reg708 <= reg641[(4'h8):(1'h1)];
            end
          else
            begin
              reg708 <= $signed(reg649);
              reg709 = ($unsigned(reg649) && $unsigned(reg686[(1'h1):(1'h0)]));
              reg710 <= $unsigned($unsigned((7'h45)));
              reg711 <= reg668[(5'h12):(5'h10)];
            end
          for (forvar712 = (1'h0); (forvar712 < (2'h2)); forvar712 = (forvar712 + (1'h1)))
            begin
              reg713 = ($signed(reg684) >= ($signed($unsigned(reg634[(2'h2):(1'h1)])) == ({reg705,
                  reg623} == reg682[(5'h13):(4'h8)])));
              reg714 = (reg645[(1'h1):(1'h1)] ?
                  (((reg675 ^ $unsigned(reg689)) ?
                          (reg634 + (reg590 > reg683)) : ({reg704,
                              wire702} >>> reg683[(2'h3):(1'h0)])) ?
                      $unsigned(wire618) : $unsigned(((!wire702) * $signed(wire617)))) : wire701);
              reg715 <= ($unsigned((|({(8'hbd), reg642} ?
                  ((7'h49) ?
                      reg596 : reg697) : reg699[(4'h9):(3'h7)]))) > $unsigned(reg613));
            end
        end
      reg716 <= $unsigned((({(~|(8'haf)), $unsigned((7'h41))} ?
          ((wire701 ? reg714 : reg612) ?
              $signed(reg594) : wire583) : reg645[(1'h1):(1'h1)]) < ((!(&(8'hb0))) - ((~reg654) ?
          $signed(forvar703) : wire579[(3'h5):(1'h0)]))));
      reg717 <= (7'h44);
      for (forvar718 = (1'h0); (forvar718 < (3'h4)); forvar718 = (forvar718 + (1'h1)))
        begin
          reg719 = ((~{$signed($signed((8'ha9)))}) ?
              reg623[(4'hc):(4'hc)] : (8'hb6));
          if ($signed(reg660))
            begin
              reg720 = {($signed({$signed(reg630),
                      reg669}) & (($signed(wire580) | reg632[(3'h5):(3'h5)]) != (-(-wire591))))};
              reg721 = (-$signed((reg710[(3'h6):(1'h1)] << (|reg586))));
              reg722 = reg704;
            end
          else
            begin
              reg723 <= $signed(((($unsigned(reg631) & $signed(reg698)) ?
                      ((8'hb0) <<< ((8'hbd) >>> reg607)) : $unsigned($unsigned(reg686))) ?
                  ((^~((8'ha3) || (8'hb7))) || $signed(((8'haf) & reg719))) : reg710[(4'ha):(1'h0)]));
              reg724 <= $unsigned($unsigned(reg709[(4'h8):(3'h6)]));
              reg725 <= ((({{(8'ha7), reg698}, $unsigned(wire648)} ?
                          ($unsigned(reg698) == (|reg708)) : reg683) ?
                      $unsigned(reg724[(2'h3):(1'h0)]) : (reg629[(2'h3):(2'h2)] ?
                          (~|$signed(wire591)) : ((~reg669) ?
                              reg719 : (reg722 > reg613)))) ?
                  ({$signed((8'ha7)),
                          ($signed(reg637) ? (wire580 >= reg682) : {reg671})} ?
                      ((8'hae) ? {wire579} : wire618) : {($signed((8'hac)) ?
                              $signed(forvar703) : $signed((8'ha3))),
                          reg634[(3'h4):(2'h3)]}) : (reg593 ?
                      (~reg697[(1'h1):(1'h0)]) : reg649));
              reg726 = reg641;
              reg727 = (!(wire585[(3'h5):(3'h4)] <<< $signed(((reg612 ?
                  forvar718 : reg723) && reg645))));
            end
          if ($signed(reg724[(4'he):(3'h5)]))
            begin
              reg728 = ($unsigned(reg664[(3'h5):(3'h4)]) ?
                  $unsigned((~&$unsigned((reg602 || reg723)))) : reg720[(2'h2):(1'h0)]);
              reg729 <= $unsigned((^~((+(reg713 <= reg705)) ?
                  (!reg602[(3'h5):(2'h2)]) : ((reg668 ? reg614 : reg670) ?
                      $signed(reg721) : (reg671 * reg686)))));
              reg730 = $unsigned((reg706 >>> $unsigned(($signed(reg669) ?
                  (reg719 - reg646) : reg654))));
              reg731 = (+(~^(&$unsigned(reg717[(3'h6):(3'h4)]))));
            end
          else
            begin
              reg728 = (reg634[(1'h0):(1'h0)] ?
                  reg645[(2'h3):(2'h3)] : $signed($signed($unsigned({reg641}))));
              reg730 = $signed(($unsigned(($unsigned(wire617) == (+wire584))) <= forvar703));
              reg732 <= ($unsigned(forvar712[(4'ha):(4'h9)]) ?
                  $signed((~($signed(reg649) <<< (|reg616)))) : (($signed(forvar718) * (&$unsigned(reg631))) ?
                      wire581 : (|reg719)));
              reg733 <= ({reg689[(3'h4):(2'h2)], $signed((~^reg641))} ?
                  ({$signed((reg683 >>> reg590)), (|(~^reg669))} ?
                      reg593 : reg593) : (wire701[(2'h3):(2'h3)] ?
                      reg726[(4'h8):(1'h0)] : reg616[(3'h5):(1'h0)]));
            end
        end
    end
  assign wire734 = reg724[(3'h7):(1'h0)];
  assign wire735 = $unsigned(reg671[(3'h4):(3'h4)]);
  assign wire736 = $signed($unsigned(wire585[(1'h0):(1'h0)]));
endmodule