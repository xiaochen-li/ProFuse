(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param1172 = {((({(8'hb8), (8'hba)} ? (~(8'hb6)) : ((8'hbd) ? (8'haa) : (8'haf))) <<< ((^(7'h40)) >>> ((8'hba) ? (8'had) : (8'hb7)))) ? ({((8'hb9) ? (8'ha8) : (8'hb9)), ((8'hbb) - (8'hb1))} ? (((8'ha9) - (8'hb1)) ? ((8'h9d) ? (8'ha1) : (8'hb1)) : (+(8'h9c))) : (~|((8'hbc) < (8'h9f)))) : ((+(~(8'hb0))) ? {(8'h9d)} : (|(~^(8'hba))))), (-{(((7'h40) == (8'haf)) ? {(8'ha6)} : (^(8'hbd)))})} )
(y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h518):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire4;
  input wire [(5'h15):(1'h0)] wire3;
  input wire signed [(4'hf):(1'h0)] wire2;
  input wire signed [(4'hb):(1'h0)] wire1;
  input wire signed [(5'h14):(1'h0)] wire0;
  wire signed [(5'h15):(1'h0)] wire1171;
  wire [(4'hd):(1'h0)] wire1169;
  reg signed [(3'h4):(1'h0)] reg1168 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1167 = (1'h0);
  reg [(3'h7):(1'h0)] reg1166 = (1'h0);
  reg [(5'h11):(1'h0)] reg1165 = (1'h0);
  reg [(5'h10):(1'h0)] reg1164 = (1'h0);
  reg [(3'h6):(1'h0)] reg1163 = (1'h0);
  wire [(5'h11):(1'h0)] wire1162;
  wire signed [(4'he):(1'h0)] wire1161;
  wire signed [(4'hc):(1'h0)] wire1159;
  reg [(3'h7):(1'h0)] reg1158 = (1'h0);
  reg [(4'hb):(1'h0)] reg1157 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1156 = (1'h0);
  reg [(4'hb):(1'h0)] reg1155 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1154 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1153 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1152 = (1'h0);
  reg [(4'h9):(1'h0)] reg1151 = (1'h0);
  reg [(5'h10):(1'h0)] reg1150 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1149 = (1'h0);
  reg [(5'h13):(1'h0)] reg1148 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1147 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1146 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1145 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1144 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1143 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1142 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1141 = (1'h0);
  wire signed [(4'hc):(1'h0)] wire1139;
  reg [(3'h5):(1'h0)] reg499 = (1'h0);
  reg [(5'h11):(1'h0)] reg498 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg497 = (1'h0);
  reg [(4'hc):(1'h0)] reg496 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg495 = (1'h0);
  wire signed [(4'ha):(1'h0)] wire494;
  wire [(4'he):(1'h0)] wire492;
  reg [(4'h8):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg71 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg70 = (1'h0);
  reg [(4'hf):(1'h0)] reg69 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg68 = (1'h0);
  reg [(2'h3):(1'h0)] forvar67 = (1'h0);
  reg [(2'h2):(1'h0)] reg66 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar65 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg64 = (1'h0);
  reg [(4'ha):(1'h0)] reg63 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar62 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg61 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire60;
  reg [(4'hc):(1'h0)] reg55 = (1'h0);
  reg [(4'hd):(1'h0)] reg49 = (1'h0);
  reg [(5'h13):(1'h0)] reg47 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar45 = (1'h0);
  reg [(2'h2):(1'h0)] reg59 = (1'h0);
  reg [(5'h12):(1'h0)] reg58 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg57 = (1'h0);
  reg [(4'h8):(1'h0)] reg56 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar55 = (1'h0);
  reg [(4'hd):(1'h0)] reg54 = (1'h0);
  reg [(4'h8):(1'h0)] reg53 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg52 = (1'h0);
  reg [(3'h4):(1'h0)] reg51 = (1'h0);
  reg [(4'hb):(1'h0)] reg50 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar49 = (1'h0);
  reg [(2'h3):(1'h0)] reg48 = (1'h0);
  reg [(2'h2):(1'h0)] forvar47 = (1'h0);
  reg [(3'h5):(1'h0)] reg46 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg45 = (1'h0);
  reg [(4'h8):(1'h0)] reg44 = (1'h0);
  reg [(5'h15):(1'h0)] reg43 = (1'h0);
  reg [(5'h15):(1'h0)] reg42 = (1'h0);
  reg [(4'hc):(1'h0)] reg41 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar40 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar39 = (1'h0);
  reg [(4'hd):(1'h0)] reg38 = (1'h0);
  reg [(4'hf):(1'h0)] reg37 = (1'h0);
  reg [(2'h2):(1'h0)] reg36 = (1'h0);
  reg [(5'h14):(1'h0)] reg35 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg34 = (1'h0);
  reg [(5'h15):(1'h0)] reg33 = (1'h0);
  reg [(3'h5):(1'h0)] reg32 = (1'h0);
  reg [(5'h11):(1'h0)] reg31 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg30 = (1'h0);
  reg [(4'h9):(1'h0)] forvar29 = (1'h0);
  reg [(4'hf):(1'h0)] forvar28 = (1'h0);
  reg [(5'h11):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg26 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar25 = (1'h0);
  reg [(5'h11):(1'h0)] reg24 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg23 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg22 = (1'h0);
  reg [(5'h10):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg19 = (1'h0);
  reg [(4'hf):(1'h0)] reg18 = (1'h0);
  reg [(4'hc):(1'h0)] reg17 = (1'h0);
  reg [(3'h7):(1'h0)] reg16 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg15 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar14 = (1'h0);
  reg [(5'h14):(1'h0)] reg13 = (1'h0);
  reg [(5'h10):(1'h0)] forvar12 = (1'h0);
  reg [(4'hd):(1'h0)] reg11 = (1'h0);
  reg [(4'he):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg9 = (1'h0);
  reg [(5'h13):(1'h0)] reg8 = (1'h0);
  reg [(4'he):(1'h0)] forvar7 = (1'h0);
  reg [(2'h3):(1'h0)] forvar6 = (1'h0);
  wire [(5'h11):(1'h0)] wire5;
  assign y = {wire1171,
                 wire1169,
                 reg1168,
                 reg1167,
                 reg1166,
                 reg1165,
                 reg1164,
                 reg1163,
                 wire1162,
                 wire1161,
                 wire1159,
                 reg1158,
                 reg1157,
                 reg1156,
                 reg1155,
                 reg1154,
                 forvar1153,
                 forvar1152,
                 reg1151,
                 reg1150,
                 reg1149,
                 reg1148,
                 reg1147,
                 reg1146,
                 forvar1145,
                 reg1144,
                 reg1143,
                 forvar1142,
                 forvar1141,
                 wire1139,
                 reg499,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 wire494,
                 wire492,
                 reg65,
                 reg72,
                 reg71,
                 reg70,
                 reg69,
                 reg68,
                 forvar67,
                 reg66,
                 forvar65,
                 reg64,
                 reg63,
                 forvar62,
                 reg61,
                 wire60,
                 reg55,
                 reg49,
                 reg47,
                 forvar45,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 forvar55,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 forvar49,
                 reg48,
                 forvar47,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 forvar40,
                 forvar39,
                 reg38,
                 reg37,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 forvar29,
                 forvar28,
                 reg27,
                 reg26,
                 forvar25,
                 reg24,
                 reg23,
                 reg22,
                 reg21,
                 reg20,
                 reg19,
                 reg18,
                 reg17,
                 reg16,
                 reg15,
                 forvar14,
                 reg13,
                 forvar12,
                 reg11,
                 reg10,
                 reg9,
                 reg8,
                 forvar7,
                 forvar6,
                 wire5,
                 (1'h0)};
  assign wire5 = (wire1 ?
                     wire1 : $signed(({$signed(wire4)} ^ (^~$unsigned(wire0)))));
  always
    @(posedge clk) begin
      for (forvar6 = (1'h0); (forvar6 < (1'h0)); forvar6 = (forvar6 + (1'h1)))
        begin
          for (forvar7 = (1'h0); (forvar7 < (2'h3)); forvar7 = (forvar7 + (1'h1)))
            begin
              reg8 = (|$unsigned($unsigned(($unsigned(wire3) > (^~wire0)))));
              reg9 <= ($signed((~({(8'ha7)} ? forvar6 : (^reg8)))) ?
                  {(8'hbb), wire2} : $unsigned("kp91tMW9KP19kr"));
              reg10 <= forvar6[(1'h0):(1'h0)];
              reg11 <= ($unsigned((|forvar7)) ?
                  (-reg10[(3'h6):(2'h3)]) : forvar6);
            end
        end
      for (forvar12 = (1'h0); (forvar12 < (3'h4)); forvar12 = (forvar12 + (1'h1)))
        begin
          reg13 <= $unsigned({((~|"4qyTHLyIy1YuvN9zIIH") ?
                  {$unsigned(reg8)} : {$signed((8'hbb))})});
          for (forvar14 = (1'h0); (forvar14 < (1'h1)); forvar14 = (forvar14 + (1'h1)))
            begin
              reg15 <= ({$unsigned($signed($unsigned(forvar6)))} ?
                  ($unsigned(wire2[(4'hc):(4'hc)]) ?
                      ($unsigned($unsigned(reg13)) ?
                          (~reg13) : $unsigned({wire4,
                              forvar6})) : wire0) : $unsigned({$signed($signed(wire0)),
                      ((forvar7 ? wire4 : forvar7) ?
                          forvar6[(1'h1):(1'h0)] : forvar6[(1'h0):(1'h0)])}));
              reg16 <= (8'ha8);
              reg17 = (!$unsigned($unsigned(reg11[(3'h5):(1'h0)])));
              reg18 = (wire2[(4'hb):(1'h0)] ?
                  (8'hb1) : $signed(({{wire2, reg8}, (wire4 < wire5)} ?
                      $signed(((8'haf) ?
                          wire3 : forvar6)) : reg9[(3'h7):(2'h3)])));
            end
          if ((((-wire4) == $signed(wire4)) >= $unsigned((($signed(reg15) != (~|(8'hbf))) ?
              ("kbMw3a5U3" ? {reg17} : "9KM") : ((^wire2) ?
                  $unsigned(reg9) : wire4)))))
            begin
              reg19 <= ((~&(reg8 ?
                  (~^$unsigned(wire3)) : wire4)) - reg15[(3'h4):(1'h0)]);
              reg20 = ($unsigned(($signed((reg11 >= wire5)) ?
                  (~&(+wire3)) : forvar12[(3'h7):(3'h6)])) >> reg16[(3'h6):(3'h5)]);
              reg21 = (~|$signed($signed((forvar6 <= $unsigned(wire2)))));
              reg22 <= reg11[(2'h3):(1'h0)];
              reg23 = reg18;
            end
          else
            begin
              reg19 <= {((~^{{reg11}}) ?
                      forvar6[(2'h3):(1'h0)] : ((^(!(8'haa))) + (&(reg13 ?
                          forvar12 : reg10)))),
                  (+reg20)};
              reg20 <= reg20[(2'h3):(2'h2)];
            end
          reg24 = $unsigned($unsigned("tpnISFFFUTKllBZa"));
          for (forvar25 = (1'h0); (forvar25 < (1'h1)); forvar25 = (forvar25 + (1'h1)))
            begin
              reg26 <= $signed(((reg21[(3'h7):(3'h5)] ?
                      $unsigned((reg16 ? wire0 : wire1)) : "Ksyim2Yu") ?
                  forvar14 : reg24[(4'hd):(3'h5)]));
              reg27 <= wire2;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar28 = (1'h0); (forvar28 < (1'h1)); forvar28 = (forvar28 + (1'h1)))
        begin
          for (forvar29 = (1'h0); (forvar29 < (2'h3)); forvar29 = (forvar29 + (1'h1)))
            begin
              reg30 = (wire4 ?
                  (-forvar6[(1'h0):(1'h0)]) : reg18[(4'he):(4'hc)]);
              reg31 <= ((8'had) <<< $signed(forvar7));
              reg32 <= {{$signed({forvar12[(4'hb):(4'ha)]}),
                      (reg22 ?
                          $signed(forvar25[(3'h5):(1'h1)]) : (wire1 <<< (forvar14 - wire2)))},
                  (wire0[(2'h3):(1'h1)] ^~ $signed($signed((reg26 || forvar14))))};
            end
          reg33 = ((wire1 ?
              forvar25[(3'h4):(2'h3)] : (($unsigned(reg21) ?
                      $signed(reg15) : reg15) ?
                  reg9[(2'h2):(1'h1)] : $unsigned((!wire1)))) == $signed({((-(8'ha0)) ?
                  $unsigned(forvar14) : reg17[(2'h3):(1'h0)])}));
          reg34 <= $unsigned(reg24);
          reg35 <= $unsigned($unsigned((reg13[(4'hb):(1'h1)] || (-(forvar25 & wire1)))));
          if ((wire0 ?
              $unsigned(forvar14) : (((!reg33[(4'hb):(4'hb)]) ?
                      (!reg21[(4'hc):(1'h1)]) : $signed((forvar14 ?
                          forvar29 : reg22))) ?
                  $signed(((^(7'h43)) ?
                      {reg22,
                          reg11} : $signed((8'ha9)))) : (!(reg15[(3'h5):(2'h3)] ^~ {reg23,
                      wire4})))))
            begin
              reg36 = $unsigned((8'haf));
              reg37 <= forvar14[(2'h3):(2'h2)];
              reg38 = $signed((({(reg8 != reg15)} ?
                      (~^$unsigned(reg35)) : {(~reg10),
                          ((8'ha4) ? reg34 : reg36)}) ?
                  reg24 : (~&$signed($unsigned((8'hb7))))));
            end
          else
            begin
              reg36 <= ((|(reg31[(3'h7):(3'h5)] ?
                  $unsigned(reg18) : reg13)) | $signed(($unsigned((reg35 ?
                  forvar29 : reg19)) > (8'hab))));
              reg37 <= wire4;
            end
        end
      for (forvar39 = (1'h0); (forvar39 < (2'h3)); forvar39 = (forvar39 + (1'h1)))
        begin
          for (forvar40 = (1'h0); (forvar40 < (1'h0)); forvar40 = (forvar40 + (1'h1)))
            begin
              reg41 = (~&($unsigned(($signed(forvar12) >>> reg36[(2'h2):(2'h2)])) ?
                  (~&(^~$unsigned(reg34))) : (reg13[(5'h13):(3'h5)] >> (!$signed(reg23)))));
            end
          if (((^~$unsigned((+"3EAYiLm2sZs"))) ? reg19 : reg35))
            begin
              reg42 <= "SYyAAtyZLR46";
              reg43 <= (~|$unsigned(reg9));
              reg44 <= $signed(forvar39[(3'h4):(3'h4)]);
            end
          else
            begin
              reg42 <= $signed($signed((reg33 - {{forvar39, wire0}})));
            end
        end
      if ((~|reg23))
        begin
          reg45 = $unsigned(reg27[(4'hb):(2'h3)]);
          reg46 = $unsigned((^wire3));
          for (forvar47 = (1'h0); (forvar47 < (2'h2)); forvar47 = (forvar47 + (1'h1)))
            begin
              reg48 <= $unsigned({reg43[(4'ha):(2'h3)]});
            end
          for (forvar49 = (1'h0); (forvar49 < (2'h3)); forvar49 = (forvar49 + (1'h1)))
            begin
              reg50 = ({reg38, $signed(forvar39)} ?
                  reg26 : (wire4[(1'h0):(1'h0)] & wire1));
              reg51 <= $unsigned(($unsigned(reg26) <= $signed(((forvar29 ?
                  forvar49 : reg9) & (^(8'h9e))))));
              reg52 <= ($unsigned($signed((&$signed(reg50)))) ^~ "7tSY");
              reg53 <= (~&$unsigned($signed($unsigned($signed(forvar14)))));
              reg54 = $unsigned($signed(reg22));
            end
          for (forvar55 = (1'h0); (forvar55 < (2'h2)); forvar55 = (forvar55 + (1'h1)))
            begin
              reg56 <= {reg48[(2'h2):(1'h1)]};
              reg57 = reg15;
              reg58 <= $unsigned(forvar40);
              reg59 <= (8'ha4);
            end
        end
      else
        begin
          for (forvar45 = (1'h0); (forvar45 < (1'h1)); forvar45 = (forvar45 + (1'h1)))
            begin
              reg46 = ((^reg17) >>> ((^~wire5[(4'ha):(2'h3)]) ~^ $unsigned(((-forvar49) > reg31))));
              reg47 <= forvar28;
              reg48 <= wire0[(3'h5):(2'h3)];
              reg49 = (~$unsigned(reg13));
              reg50 <= reg10;
            end
          reg51 <= reg32;
          reg52 = (reg9 ~^ $signed((($unsigned(reg58) && ((7'h41) ?
              (8'hb2) : reg47)) ~^ {forvar40[(2'h2):(1'h0)]})));
          if ((~|((reg30[(2'h2):(1'h1)] + forvar14) ?
              $unsigned((8'hbd)) : {(!$signed(reg50))})))
            begin
              reg53 <= ($signed("FSd2dshhWYcU") != (8'ha1));
              reg54 <= (^~(~(reg16 ? $signed((^~reg37)) : "WZT0VyV9OY8Lz2tl")));
              reg55 = forvar40[(4'h9):(4'h8)];
              reg56 = (("NCGCcwXvMmV3DdMZRbYO" ?
                      (reg55[(4'hc):(2'h3)] ^ (reg30[(4'h8):(3'h5)] >= reg42[(4'hc):(4'h8)])) : ((8'h9f) ?
                          $unsigned($signed(reg43)) : $signed((~forvar49)))) ?
                  reg48[(1'h1):(1'h1)] : (reg34[(3'h4):(2'h2)] ?
                      $signed({$signed(reg38),
                          (reg49 ^ reg11)}) : $signed((reg58[(4'hf):(1'h0)] ?
                          (!forvar29) : (^forvar45)))));
              reg57 = (8'h9e);
            end
          else
            begin
              reg53 = wire4;
              reg54 = ($signed(((|reg32) ? (8'hb0) : {(+reg46)})) ?
                  reg36[(1'h0):(1'h0)] : (forvar29 << {$signed(reg23),
                      $signed((reg16 ? reg52 : reg58))}));
              reg55 <= $unsigned(reg11);
            end
        end
    end
  assign wire60 = forvar12;
  always
    @(posedge clk) begin
      if (((^{(-forvar39[(2'h3):(1'h1)]),
          ($signed(reg38) ?
              $signed(reg50) : (wire3 > forvar49))}) != (!wire0[(5'h13):(4'hc)])))
        begin
          reg61 <= $unsigned(reg11);
          for (forvar62 = (1'h0); (forvar62 < (2'h2)); forvar62 = (forvar62 + (1'h1)))
            begin
              reg63 <= $signed(($unsigned(reg18[(4'h9):(1'h0)]) >> $unsigned(reg23[(1'h0):(1'h0)])));
            end
          reg64 = $unsigned(reg31[(3'h7):(3'h5)]);
          for (forvar65 = (1'h0); (forvar65 < (2'h2)); forvar65 = (forvar65 + (1'h1)))
            begin
              reg66 <= (reg23[(3'h5):(1'h0)] ? reg47 : "msnfRTSWdmwTtfZJKOl");
            end
          for (forvar67 = (1'h0); (forvar67 < (2'h3)); forvar67 = (forvar67 + (1'h1)))
            begin
              reg68 <= $unsigned({(reg32[(2'h3):(1'h0)] ?
                      (^~reg52[(1'h1):(1'h1)]) : (wire60 - forvar14[(1'h1):(1'h0)])),
                  reg15[(2'h3):(1'h1)]});
              reg69 <= (($unsigned($unsigned((wire0 > (8'hac)))) * (($signed(forvar25) ?
                  $signed(reg63) : wire2) <= ($signed(reg33) < $unsigned(reg19)))) ^~ {reg64,
                  ($unsigned($signed((8'hb1))) ?
                      reg24[(4'h8):(1'h0)] : ((reg23 | forvar39) ?
                          forvar25 : wire3))});
              reg70 <= forvar29;
              reg71 = (($unsigned(((reg22 != reg45) ?
                      (forvar29 ? forvar12 : reg22) : {reg36,
                          reg9})) << $unsigned((reg32 ?
                      (reg36 ^ (8'hb6)) : reg58))) ?
                  $unsigned(reg70[(4'h9):(1'h0)]) : (~^($signed(reg45) ?
                      ($signed(reg11) >= forvar14[(2'h3):(1'h0)]) : (~&(reg27 && reg56)))));
              reg72 <= {($signed(({reg18} << forvar14)) > {(~reg8[(4'ha):(2'h3)])}),
                  ("LXte6N" <<< reg18)};
            end
        end
      else
        begin
          reg61 <= ((8'ha3) ?
              $signed(({$signed(forvar7),
                  $signed(reg55)} != wire1)) : ((reg26[(4'hf):(4'ha)] >> (^(&(8'hb0)))) ?
                  $unsigned($signed($unsigned(reg30))) : $unsigned((8'hb0))));
          for (forvar62 = (1'h0); (forvar62 < (2'h2)); forvar62 = (forvar62 + (1'h1)))
            begin
              reg63 <= reg55[(4'hc):(3'h7)];
              reg64 <= $unsigned((reg50[(4'h9):(1'h0)] ?
                  ($unsigned($unsigned(reg26)) < reg44[(1'h1):(1'h1)]) : reg42[(4'h9):(2'h3)]));
            end
          reg65 = $unsigned((&$signed({$unsigned(reg16)})));
          reg66 = reg9[(2'h2):(1'h0)];
        end
    end
  module73 modinst493 (wire492, clk, reg26, reg31, forvar12, reg44);
  assign wire494 = (($unsigned(reg32) ?
                       reg15 : {($signed(reg31) ?
                               (forvar12 ?
                                   (8'hac) : reg10) : $signed(reg45))}) == $unsigned((((+reg15) > "ao1l") >> ($unsigned(forvar14) ?
                       reg35 : forvar6[(1'h1):(1'h0)]))));
  always
    @(posedge clk) begin
      reg495 <= reg65[(3'h5):(2'h2)];
      reg496 = (wire1 ?
          ((+($unsigned(reg17) > (reg56 & reg26))) ?
              (~$unsigned(((8'hb7) << forvar28))) : $signed((^$unsigned(reg64)))) : {reg59,
              $signed(reg51)});
      reg497 = {reg10};
      reg498 <= {forvar62};
      reg499 <= ((~&((reg44 ?
              (reg10 ? reg55 : reg16) : (|reg16)) + (&$unsigned(reg497)))) ?
          $unsigned((^~$unsigned(forvar67[(2'h2):(2'h2)]))) : $unsigned((($signed(reg71) ?
                  $signed(reg10) : (8'h9f)) ?
              $unsigned($unsigned(reg52)) : {(forvar25 ? reg18 : (8'had))})));
    end
  module500 modinst1140 (.wire504(forvar45), .wire502(reg11), .wire503(forvar28), .y(wire1139), .wire501(reg37), .clk(clk));
  always
    @(posedge clk) begin
      for (forvar1141 = (1'h0); (forvar1141 < (2'h3)); forvar1141 = (forvar1141 + (1'h1)))
        begin
          for (forvar1142 = (1'h0); (forvar1142 < (1'h0)); forvar1142 = (forvar1142 + (1'h1)))
            begin
              reg1143 <= (!reg55);
              reg1144 <= reg55;
            end
          for (forvar1145 = (1'h0); (forvar1145 < (3'h4)); forvar1145 = (forvar1145 + (1'h1)))
            begin
              reg1146 <= ((reg53[(2'h2):(1'h1)] ?
                      {$signed((reg53 | reg11))} : {(^~$unsigned((8'hb9)))}) ?
                  forvar1145[(1'h1):(1'h0)] : reg22);
              reg1147 = (~$unsigned(((!forvar7) * {(reg44 != (8'hab))})));
              reg1148 = $signed(((({(7'h40)} - wire0) ?
                  $signed($unsigned((8'hac))) : (forvar47[(2'h2):(2'h2)] * $unsigned(reg22))) + $signed(reg497)));
              reg1149 <= forvar39[(4'hc):(3'h5)];
              reg1150 <= {{wire492,
                      ($unsigned((reg1147 & reg43)) & $signed($unsigned(forvar45)))},
                  (~&({(reg46 ? reg63 : reg10)} ?
                      (~(reg21 >> reg22)) : {reg1147, forvar12}))};
            end
          reg1151 = reg48[(2'h2):(1'h1)];
        end
      for (forvar1152 = (1'h0); (forvar1152 < (1'h0)); forvar1152 = (forvar1152 + (1'h1)))
        begin
          for (forvar1153 = (1'h0); (forvar1153 < (1'h0)); forvar1153 = (forvar1153 + (1'h1)))
            begin
              reg1154 <= $unsigned(reg61[(4'hb):(2'h3)]);
              reg1155 = forvar29[(4'h9):(4'h9)];
              reg1156 <= $signed(reg69);
              reg1157 = {(8'hab), (&$unsigned($unsigned((^~reg22))))};
              reg1158 <= $unsigned({(^~(forvar40 + (reg10 < reg46))),
                  $unsigned(($signed((8'hae)) <= (^~reg13)))});
            end
        end
    end
  module313 modinst1160 (.wire314(forvar7), .y(wire1159), .clk(clk), .wire317(forvar40), .wire316(reg22), .wire315(reg19));
  assign wire1161 = ($unsigned((forvar28 < $unsigned((wire1159 + reg1157)))) ?
                        wire0 : $signed($signed($signed((reg64 == forvar65)))));
  assign wire1162 = $signed($signed((7'h44)));
  always
    @(posedge clk) begin
      if ((-(+"wIJkTlkGMzgu6r")))
        begin
          reg1163 <= (7'h44);
          if ($unsigned({(8'h9f), (!$signed((reg495 ? reg1144 : reg63)))}))
            begin
              reg1164 <= $signed(reg10[(4'h9):(1'h0)]);
              reg1165 = reg1151[(2'h3):(1'h0)];
              reg1166 <= reg68;
              reg1167 <= $unsigned((!reg1163));
            end
          else
            begin
              reg1164 <= (reg71[(3'h7):(2'h3)] ? reg15 : {reg1156});
              reg1165 <= ({$unsigned(wire1159),
                  wire3} && reg1148[(4'hc):(1'h0)]);
              reg1166 <= ($signed(forvar12[(2'h2):(1'h1)]) >> $unsigned($signed(("dzW" - (&(8'ha8))))));
              reg1167 <= ($unsigned({$unsigned(reg16[(1'h1):(1'h1)])}) ?
                  $unsigned(forvar7) : $unsigned("uEutCneQE6fwRCJ0TA"));
            end
        end
      else
        begin
          if ((+reg33[(4'hf):(4'hf)]))
            begin
              reg1163 <= (!$unsigned(($signed($signed(reg1148)) ?
                  $unsigned("yBTWo") : reg46[(2'h2):(2'h2)])));
              reg1164 = (8'h9c);
              reg1165 <= {($signed(reg1146[(3'h6):(2'h3)]) ?
                      forvar65 : (^~$signed((forvar1142 > reg1156)))),
                  ((~|$signed((reg49 ? (8'hbc) : reg499))) ?
                      {$signed("4AVYDPcLt"),
                          $signed($signed(wire494))} : (wire1139[(3'h5):(3'h5)] ?
                          ({reg15} <<< wire492) : reg10[(3'h6):(3'h4)]))};
            end
          else
            begin
              reg1163 <= forvar6[(1'h1):(1'h1)];
              reg1164 <= (~forvar62[(4'hc):(2'h3)]);
              reg1165 <= (&(!(((reg1158 >= forvar1141) >>> (reg59 || forvar49)) <= reg1166)));
            end
        end
      reg1168 <= (8'hb9);
    end
  module73 modinst1170 (.wire74(wire1159), .y(wire1169), .wire77(reg19), .wire76(reg41), .wire75(wire492), .clk(clk));
  assign wire1171 = $unsigned("XfD");
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module500
#( parameter param1137 = ((8'had) || (^~(((~&(8'h9f)) >>> ((8'h9c) || (8'hbd))) != ((~(8'h9e)) ? {(8'h9c), (7'h40)} : (+(8'ha5))))))
, parameter param1138 = (!param1137) )
(y, clk, wire504, wire503, wire502, wire501);
  output wire [(32'h464):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire504;
  input wire signed [(4'hf):(1'h0)] wire503;
  input wire signed [(4'hd):(1'h0)] wire502;
  input wire signed [(4'hf):(1'h0)] wire501;
  wire [(2'h2):(1'h0)] wire1136;
  wire signed [(5'h15):(1'h0)] wire642;
  wire signed [(4'h8):(1'h0)] wire509;
  wire signed [(5'h10):(1'h0)] wire508;
  reg [(3'h7):(1'h0)] reg507 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg506 = (1'h0);
  reg [(5'h15):(1'h0)] reg505 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire745;
  reg signed [(4'h8):(1'h0)] forvar747 = (1'h0);
  reg [(5'h15):(1'h0)] reg748 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar749 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg750 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg751 = (1'h0);
  reg [(4'h9):(1'h0)] reg752 = (1'h0);
  reg [(3'h4):(1'h0)] reg753 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg754 = (1'h0);
  reg [(2'h3):(1'h0)] reg755 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg756 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg757 = (1'h0);
  reg [(5'h12):(1'h0)] reg758 = (1'h0);
  reg [(4'he):(1'h0)] reg759 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg760 = (1'h0);
  reg signed [(4'he):(1'h0)] reg761 = (1'h0);
  reg [(5'h11):(1'h0)] reg762 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg763 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg764 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar765 = (1'h0);
  reg [(5'h11):(1'h0)] reg766 = (1'h0);
  reg [(4'ha):(1'h0)] reg767 = (1'h0);
  reg [(2'h3):(1'h0)] forvar752 = (1'h0);
  reg [(4'ha):(1'h0)] forvar759 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar761 = (1'h0);
  reg [(5'h11):(1'h0)] reg765 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar768 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg769 = (1'h0);
  reg [(5'h13):(1'h0)] reg770 = (1'h0);
  reg [(5'h14):(1'h0)] reg771 = (1'h0);
  reg [(4'hf):(1'h0)] reg772 = (1'h0);
  reg [(5'h13):(1'h0)] forvar773 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg774 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar772 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg773 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg775 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg776 = (1'h0);
  reg [(3'h5):(1'h0)] reg777 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg778 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg779 = (1'h0);
  reg [(3'h6):(1'h0)] reg780 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire781;
  reg [(4'h9):(1'h0)] reg782 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg783 = (1'h0);
  reg [(4'ha):(1'h0)] reg784 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar785 = (1'h0);
  reg [(3'h5):(1'h0)] reg786 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg787 = (1'h0);
  reg [(4'hc):(1'h0)] reg788 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg789 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar790 = (1'h0);
  reg [(5'h14):(1'h0)] forvar791 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg792 = (1'h0);
  reg [(3'h6):(1'h0)] reg793 = (1'h0);
  reg [(4'h8):(1'h0)] reg794 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg795 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar796 = (1'h0);
  reg [(3'h7):(1'h0)] reg797 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg798 = (1'h0);
  reg [(5'h12):(1'h0)] reg799 = (1'h0);
  reg [(3'h7):(1'h0)] reg800 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg801 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg802 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar803 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg804 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg805 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg806 = (1'h0);
  reg [(4'ha):(1'h0)] reg807 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar808 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg809 = (1'h0);
  reg [(2'h3):(1'h0)] reg810 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg811 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar812 = (1'h0);
  reg [(4'hf):(1'h0)] reg813 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar814 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg815 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg816 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire817;
  wire signed [(4'hf):(1'h0)] wire999;
  wire [(5'h14):(1'h0)] wire1001;
  wire [(5'h12):(1'h0)] wire1002;
  wire [(5'h15):(1'h0)] wire1134;
  assign y = {wire1136,
                 wire642,
                 wire509,
                 wire508,
                 reg507,
                 reg506,
                 reg505,
                 wire745,
                 forvar747,
                 reg748,
                 forvar749,
                 reg750,
                 reg751,
                 reg752,
                 reg753,
                 reg754,
                 reg755,
                 reg756,
                 reg757,
                 reg758,
                 reg759,
                 reg760,
                 reg761,
                 reg762,
                 reg763,
                 reg764,
                 forvar765,
                 reg766,
                 reg767,
                 forvar752,
                 forvar759,
                 forvar761,
                 reg765,
                 forvar768,
                 reg769,
                 reg770,
                 reg771,
                 reg772,
                 forvar773,
                 reg774,
                 forvar772,
                 reg773,
                 reg775,
                 reg776,
                 reg777,
                 reg778,
                 reg779,
                 reg780,
                 wire781,
                 reg782,
                 reg783,
                 reg784,
                 forvar785,
                 reg786,
                 reg787,
                 reg788,
                 reg789,
                 forvar790,
                 forvar791,
                 reg792,
                 reg793,
                 reg794,
                 reg795,
                 forvar796,
                 reg797,
                 reg798,
                 reg799,
                 reg800,
                 reg801,
                 reg802,
                 forvar803,
                 reg804,
                 reg805,
                 reg806,
                 reg807,
                 forvar808,
                 reg809,
                 reg810,
                 reg811,
                 forvar812,
                 reg813,
                 forvar814,
                 reg815,
                 reg816,
                 wire817,
                 wire999,
                 wire1001,
                 wire1002,
                 wire1134,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg505 <= (($signed({(wire501 > wire502), (!wire502)}) ?
          wire503 : ((&wire501[(4'h9):(3'h7)]) ?
              {wire503[(1'h0):(1'h0)],
                  (wire501 ~^ wire502)} : wire503)) < {$signed(({wire502,
                  wire502} ?
              (wire501 + wire502) : (+wire502)))});
      reg506 <= $signed(reg505);
      reg507 <= reg506;
    end
  assign wire508 = wire503;
  assign wire509 = $unsigned($signed($signed($unsigned({(8'ha5), wire502}))));
  module510 modinst643 (wire642, clk, reg506, wire508, wire503, wire504, reg507);
  module644 modinst746 (.wire645(wire502), .wire646(wire504), .wire648(reg506), .y(wire745), .wire647(wire508), .clk(clk));
  always
    @(posedge clk) begin
      for (forvar747 = (1'h0); (forvar747 < (1'h1)); forvar747 = (forvar747 + (1'h1)))
        begin
          reg748 <= ((8'h9c) >>> $signed(reg506));
        end
      for (forvar749 = (1'h0); (forvar749 < (1'h0)); forvar749 = (forvar749 + (1'h1)))
        begin
          reg750 <= $unsigned($signed((+$unsigned((forvar747 ?
              wire642 : (8'hb4))))));
        end
      reg751 <= wire642;
      if ((~$unsigned((8'hbb))))
        begin
          if (wire642)
            begin
              reg752 = $unsigned(wire502);
              reg753 = (~((&$signed((wire501 <<< reg505))) ?
                  $signed($signed(reg748[(5'h11):(5'h10)])) : ((~$unsigned(reg748)) || {$unsigned(reg752)})));
              reg754 <= ((8'hb7) == forvar749[(4'hb):(1'h1)]);
            end
          else
            begin
              reg752 = ((8'ha2) >> (|(((wire745 ?
                      (8'hac) : (8'h9f)) == $unsigned(wire501)) ?
                  forvar747 : wire502)));
              reg753 = (8'ha9);
              reg754 = wire745;
            end
          if ($unsigned(($signed((^~wire642[(3'h4):(1'h0)])) - (~|$signed((reg748 < reg751))))))
            begin
              reg755 <= forvar749[(3'h7):(2'h2)];
              reg756 <= reg751;
            end
          else
            begin
              reg755 = $signed(($unsigned($unsigned("Q2AC64Ja2JnatyfbE")) ?
                  $signed($unsigned({wire503,
                      wire504})) : $signed({$signed(reg751), (+forvar749)})));
              reg756 = $signed(wire642);
              reg757 <= $unsigned((+reg506));
              reg758 <= forvar747[(2'h3):(1'h1)];
            end
          if ((wire501 ? (~&wire501) : $signed("szVo")))
            begin
              reg759 = $signed($signed(($unsigned($unsigned(reg753)) ?
                  (!(forvar747 ? reg751 : reg751)) : ((+(8'hae)) ^~ wire504))));
              reg760 = reg505[(3'h6):(1'h1)];
              reg761 = (($unsigned(reg748[(5'h12):(1'h1)]) <<< ({reg754,
                      (8'ha9)} ?
                  ($unsigned((7'h42)) ?
                      (|forvar749) : (~|reg506)) : (reg756 >= $unsigned(reg507)))) && reg757);
              reg762 = wire509;
              reg763 <= (($signed(wire504) - wire501) ~^ wire502);
            end
          else
            begin
              reg759 = wire509;
              reg760 = "U";
            end
          reg764 <= ($unsigned(((~^reg756[(1'h1):(1'h1)]) != (-(wire745 ?
                  (8'ha3) : reg758)))) ?
              $unsigned(forvar747[(3'h4):(2'h3)]) : reg505);
          for (forvar765 = (1'h0); (forvar765 < (2'h3)); forvar765 = (forvar765 + (1'h1)))
            begin
              reg766 = reg762;
              reg767 <= $unsigned($unsigned($unsigned(($signed(reg763) ?
                  ((8'had) ? reg751 : reg755) : reg753))));
            end
        end
      else
        begin
          for (forvar752 = (1'h0); (forvar752 < (1'h1)); forvar752 = (forvar752 + (1'h1)))
            begin
              reg753 <= $unsigned({{wire503[(2'h2):(2'h2)]}});
              reg754 = $unsigned(reg763);
              reg755 <= (!({"bxhK8l"} ^~ $unsigned($unsigned($unsigned(reg763)))));
              reg756 <= ($signed(reg757[(2'h2):(1'h1)]) >> "");
              reg757 <= reg767[(3'h5):(3'h5)];
            end
          reg758 <= wire745[(2'h2):(1'h0)];
          for (forvar759 = (1'h0); (forvar759 < (2'h2)); forvar759 = (forvar759 + (1'h1)))
            begin
              reg760 <= {$signed(wire502),
                  ($unsigned($unsigned($signed(reg505))) && reg759[(3'h4):(3'h4)])};
            end
          for (forvar761 = (1'h0); (forvar761 < (2'h3)); forvar761 = (forvar761 + (1'h1)))
            begin
              reg762 <= {$signed(reg762[(1'h0):(1'h0)])};
              reg763 <= reg761[(4'hd):(3'h5)];
              reg764 <= "LW0cSt5s";
              reg765 = $signed((~|((!forvar749) - (((7'h41) ?
                  reg507 : reg758) & $signed(wire745)))));
            end
          reg766 <= ($signed((reg763[(3'h7):(3'h4)] ?
              ((~reg752) - (wire509 != reg767)) : $unsigned((~reg753)))) < $unsigned(wire508[(4'he):(4'h9)]));
        end
      if (forvar749)
        begin
          for (forvar768 = (1'h0); (forvar768 < (2'h2)); forvar768 = (forvar768 + (1'h1)))
            begin
              reg769 <= (~|wire642[(4'hf):(1'h1)]);
              reg770 = reg767;
              reg771 = ((reg751[(3'h6):(2'h2)] ?
                      (|reg751[(3'h6):(1'h1)]) : ($unsigned($signed(wire642)) << $signed($unsigned(reg758)))) ?
                  forvar752 : $signed($unsigned((^~((8'hb9) < reg748)))));
              reg772 = {reg766};
            end
          for (forvar773 = (1'h0); (forvar773 < (3'h4)); forvar773 = (forvar773 + (1'h1)))
            begin
              reg774 = forvar773;
            end
        end
      else
        begin
          for (forvar768 = (1'h0); (forvar768 < (3'h4)); forvar768 = (forvar768 + (1'h1)))
            begin
              reg769 <= ({$signed({{wire508}, (reg763 >> reg764)})} ?
                  (reg760 == $unsigned(forvar761)) : $signed(((~^$unsigned(reg771)) ?
                      {$signed(reg772), $unsigned(reg769)} : "mIbt")));
              reg770 <= $unsigned(((~^forvar747) & $unsigned({(~|wire503)})));
              reg771 = reg759;
            end
          for (forvar772 = (1'h0); (forvar772 < (2'h3)); forvar772 = (forvar772 + (1'h1)))
            begin
              reg773 <= ((forvar773 != ({(reg769 ^ forvar761)} & $signed(forvar749))) ?
                  ($unsigned("l") * (~&$signed($signed(reg769)))) : (((~&(wire502 & reg507)) || ($unsigned(reg774) ?
                      (wire501 ? reg506 : wire642) : (8'ha3))) && (+reg770)));
              reg774 <= reg760;
              reg775 <= (^~((^(((8'hba) + reg772) ?
                      $unsigned(reg748) : $signed(reg755))) ?
                  ({reg760, reg764} & (forvar773[(3'h7):(3'h4)] ?
                      $signed(forvar765) : reg756)) : "m2kVnA0umHf"));
            end
          reg776 <= wire501;
          reg777 = forvar759;
          if (reg775[(4'h9):(1'h0)])
            begin
              reg778 <= reg766;
              reg779 = reg506;
              reg780 <= $unsigned((&reg758[(5'h10):(5'h10)]));
            end
          else
            begin
              reg778 <= reg772[(2'h2):(1'h1)];
              reg779 = reg760;
              reg780 <= reg506[(4'ha):(3'h5)];
            end
        end
    end
  assign wire781 = reg757[(3'h5):(1'h1)];
  always
    @(posedge clk) begin
      reg782 <= $signed((forvar768[(4'hc):(4'hc)] == ($signed((wire503 ?
              (7'h43) : reg779)) ?
          (&reg764) : (~&$signed(reg765)))));
      reg783 <= {reg755, (!{$signed({forvar752})})};
      reg784 <= (~^$unsigned(((~&(~&reg760)) && (&$unsigned(forvar773)))));
      for (forvar785 = (1'h0); (forvar785 < (2'h3)); forvar785 = (forvar785 + (1'h1)))
        begin
          if (reg779)
            begin
              reg786 = ((((reg780 ?
                      $signed((7'h44)) : forvar759[(1'h0):(1'h0)]) ?
                  reg764 : (~((8'hba) ?
                      reg775 : forvar759))) + $unsigned((!(+forvar785)))) >>> $signed($signed((reg753[(1'h1):(1'h1)] * reg774))));
              reg787 <= reg769;
              reg788 = reg770[(5'h13):(2'h2)];
              reg789 <= (-forvar768);
            end
          else
            begin
              reg786 <= reg784;
              reg787 <= reg783[(3'h4):(1'h0)];
              reg788 <= $signed(((8'hbd) ?
                  $unsigned(forvar768) : (+($signed((8'hbc)) <= (forvar772 & (8'ha0))))));
              reg789 <= $unsigned((reg766 != $unsigned($unsigned(reg759[(4'hc):(4'h8)]))));
            end
        end
      for (forvar790 = (1'h0); (forvar790 < (1'h1)); forvar790 = (forvar790 + (1'h1)))
        begin
          for (forvar791 = (1'h0); (forvar791 < (1'h1)); forvar791 = (forvar791 + (1'h1)))
            begin
              reg792 = {(|$unsigned($signed((|reg766))))};
              reg793 <= ({(reg770[(4'hc):(3'h7)] ?
                          ((~|reg784) >= ((8'hb4) ?
                              reg760 : wire503)) : ($signed(reg758) ?
                              "tn7857" : reg774[(3'h5):(1'h1)])),
                      ($signed((reg770 ?
                          reg507 : reg505)) >>> $signed($signed(reg763)))} ?
                  $unsigned((+(~^(~&reg766)))) : (($signed((+reg755)) >> (+(reg507 ?
                      wire509 : wire781))) && (^(^~$signed(reg757)))));
              reg794 <= $signed($signed((^~((forvar747 <<< reg792) ^~ (~|reg753)))));
              reg795 <= (reg752 || {$unsigned((8'hbf)), forvar752});
            end
          for (forvar796 = (1'h0); (forvar796 < (2'h3)); forvar796 = (forvar796 + (1'h1)))
            begin
              reg797 = reg759[(4'hc):(4'ha)];
              reg798 <= (reg771[(3'h7):(3'h5)] && reg756[(1'h1):(1'h0)]);
              reg799 <= $signed((~(reg769 ^~ ($unsigned((8'hbc)) & forvar747))));
              reg800 <= {reg772};
              reg801 <= $signed((&$unsigned($unsigned((+reg767)))));
            end
          reg802 = $signed((wire781 ~^ ((((8'hb4) ^~ reg756) << ((7'h43) > (8'ha7))) ?
              ($unsigned((8'hb5)) ?
                  $signed(reg800) : reg756[(4'h8):(3'h5)]) : (reg766 ?
                  reg763 : reg788))));
          for (forvar803 = (1'h0); (forvar803 < (2'h2)); forvar803 = (forvar803 + (1'h1)))
            begin
              reg804 <= reg756;
              reg805 = ({$signed({(forvar796 ? forvar785 : reg765),
                          {forvar790, forvar747}}),
                      wire642} ?
                  $signed((~^$signed(reg802[(1'h1):(1'h0)]))) : $unsigned((((reg774 >= (8'hb9)) != wire781[(1'h1):(1'h0)]) << reg763)));
            end
          reg806 <= ($signed(((wire508[(4'hb):(3'h5)] ?
                  (!reg752) : (reg798 ?
                      (8'hb1) : reg767)) && $unsigned($unsigned(wire508)))) ?
              reg783[(4'h8):(2'h3)] : reg505);
        end
    end
  always
    @(posedge clk) begin
      reg807 <= ((forvar796 ?
          $signed($signed({wire502,
              reg789})) : $unsigned(((reg802 >> wire642) ^ (forvar747 ?
              reg773 : reg761)))) != wire509[(2'h3):(1'h1)]);
      if (reg794)
        begin
          for (forvar808 = (1'h0); (forvar808 < (1'h1)); forvar808 = (forvar808 + (1'h1)))
            begin
              reg809 = ((forvar773 ^ reg793) && reg773);
              reg810 = {{(^$signed(reg776[(5'h14):(4'hd)]))}};
              reg811 <= forvar773[(4'h8):(2'h2)];
            end
        end
      else
        begin
          for (forvar808 = (1'h0); (forvar808 < (1'h1)); forvar808 = (forvar808 + (1'h1)))
            begin
              reg809 = $signed(reg804[(3'h5):(2'h2)]);
              reg810 <= $unsigned(reg752);
              reg811 <= reg806[(2'h2):(2'h2)];
            end
          for (forvar812 = (1'h0); (forvar812 < (3'h4)); forvar812 = (forvar812 + (1'h1)))
            begin
              reg813 = forvar768;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar814 = (1'h0); (forvar814 < (3'h4)); forvar814 = (forvar814 + (1'h1)))
        begin
          reg815 <= wire508[(4'h8):(3'h4)];
        end
      reg816 <= forvar790;
    end
  assign wire817 = (-reg769[(3'h5):(2'h3)]);
  module818 modinst1000 (.clk(clk), .y(wire999), .wire822(reg505), .wire821(reg767), .wire819(forvar814), .wire820(reg751));
  assign wire1001 = $unsigned((forvar765 ?
                        wire999 : ($signed("cgAyIYcRzrSKRhOdknW") ~^ (7'h40))));
  assign wire1002 = {$signed(reg779), reg794};
  module1003 modinst1135 (.clk(clk), .wire1008(reg783), .wire1006(reg799), .y(wire1134), .wire1005(reg776), .wire1004(wire509), .wire1007(reg782));
  assign wire1136 = $unsigned({(~|reg758[(4'hb):(3'h7)]),
                        ($signed((reg802 ? reg748 : forvar759)) - (-(reg751 ?
                            forvar768 : forvar796)))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module73  (y, clk, wire77, wire76, wire75, wire74);
  output wire [(32'h4e4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire77;
  input wire [(3'h5):(1'h0)] wire76;
  input wire signed [(4'he):(1'h0)] wire75;
  input wire signed [(4'h8):(1'h0)] wire74;
  wire signed [(4'hc):(1'h0)] wire491;
  wire signed [(5'h13):(1'h0)] wire490;
  wire [(3'h5):(1'h0)] wire489;
  wire [(3'h6):(1'h0)] wire488;
  wire [(4'ha):(1'h0)] wire487;
  wire [(3'h7):(1'h0)] wire486;
  wire [(3'h5):(1'h0)] wire485;
  wire signed [(5'h14):(1'h0)] wire484;
  reg signed [(2'h2):(1'h0)] reg483 = (1'h0);
  reg [(3'h5):(1'h0)] reg482 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg481 = (1'h0);
  reg [(4'he):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg479 = (1'h0);
  reg [(3'h4):(1'h0)] reg478 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg477 = (1'h0);
  reg [(3'h4):(1'h0)] forvar476 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg475 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg474 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg473 = (1'h0);
  reg [(4'hf):(1'h0)] reg472 = (1'h0);
  reg signed [(4'he):(1'h0)] reg471 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar470 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg469 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg468 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg467 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg466 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg465 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg464 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg463 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg462 = (1'h0);
  reg [(3'h5):(1'h0)] reg461 = (1'h0);
  reg [(3'h7):(1'h0)] reg460 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar459 = (1'h0);
  reg [(5'h14):(1'h0)] reg458 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar457 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg456 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg455 = (1'h0);
  reg [(3'h7):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg453 = (1'h0);
  reg [(4'hf):(1'h0)] reg452 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg451 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg450 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar449 = (1'h0);
  reg [(2'h2):(1'h0)] reg448 = (1'h0);
  reg [(3'h7):(1'h0)] reg447 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg446 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg445 = (1'h0);
  reg [(4'hc):(1'h0)] reg444 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg443 = (1'h0);
  reg [(3'h5):(1'h0)] reg442 = (1'h0);
  reg [(3'h4):(1'h0)] reg441 = (1'h0);
  reg [(4'h8):(1'h0)] forvar440 = (1'h0);
  reg [(5'h12):(1'h0)] reg439 = (1'h0);
  reg [(4'hd):(1'h0)] reg438 = (1'h0);
  reg [(3'h6):(1'h0)] reg437 = (1'h0);
  reg [(2'h2):(1'h0)] forvar436 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire434;
  wire [(4'hb):(1'h0)] wire312;
  reg [(4'hd):(1'h0)] reg311 = (1'h0);
  reg [(3'h5):(1'h0)] reg310 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg309 = (1'h0);
  reg [(3'h4):(1'h0)] reg308 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg307 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg306 = (1'h0);
  reg [(5'h12):(1'h0)] reg305 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg304 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg303 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg302 = (1'h0);
  reg [(4'ha):(1'h0)] reg301 = (1'h0);
  reg [(5'h15):(1'h0)] reg300 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg299 = (1'h0);
  reg [(4'h8):(1'h0)] forvar298 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg297 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg296 = (1'h0);
  reg [(5'h15):(1'h0)] reg295 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg294 = (1'h0);
  reg [(2'h3):(1'h0)] forvar293 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar292 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg291 = (1'h0);
  reg [(5'h14):(1'h0)] reg290 = (1'h0);
  reg [(5'h10):(1'h0)] reg289 = (1'h0);
  reg [(2'h3):(1'h0)] reg288 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg287 = (1'h0);
  reg [(4'he):(1'h0)] reg286 = (1'h0);
  reg [(2'h3):(1'h0)] reg285 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar284 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg283 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg282 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg281 = (1'h0);
  reg [(4'hb):(1'h0)] reg280 = (1'h0);
  reg [(2'h2):(1'h0)] reg279 = (1'h0);
  reg [(4'ha):(1'h0)] forvar278 = (1'h0);
  reg [(4'hb):(1'h0)] forvar277 = (1'h0);
  reg [(4'hd):(1'h0)] reg276 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg275 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg274 = (1'h0);
  reg [(4'hd):(1'h0)] reg273 = (1'h0);
  reg [(5'h12):(1'h0)] forvar272 = (1'h0);
  reg [(5'h13):(1'h0)] forvar271 = (1'h0);
  reg signed [(4'he):(1'h0)] reg270 = (1'h0);
  reg [(3'h5):(1'h0)] reg269 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg268 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg267 = (1'h0);
  reg [(4'hd):(1'h0)] reg266 = (1'h0);
  reg [(5'h10):(1'h0)] reg265 = (1'h0);
  reg [(5'h12):(1'h0)] forvar264 = (1'h0);
  reg [(5'h10):(1'h0)] reg263 = (1'h0);
  reg [(5'h13):(1'h0)] reg262 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar261 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar259 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg258 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar257 = (1'h0);
  wire signed [(5'h10):(1'h0)] wire256;
  wire signed [(4'hc):(1'h0)] wire255;
  wire signed [(3'h6):(1'h0)] wire254;
  wire signed [(5'h14):(1'h0)] wire252;
  wire signed [(4'hf):(1'h0)] wire79;
  wire [(4'he):(1'h0)] wire78;
  assign y = {wire491,
                 wire490,
                 wire489,
                 wire488,
                 wire487,
                 wire486,
                 wire485,
                 wire484,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 reg479,
                 reg478,
                 reg477,
                 forvar476,
                 reg475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 forvar470,
                 reg469,
                 reg468,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 forvar459,
                 reg458,
                 forvar457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 forvar449,
                 reg448,
                 reg447,
                 reg446,
                 reg445,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 forvar440,
                 reg439,
                 reg438,
                 reg437,
                 forvar436,
                 wire434,
                 wire312,
                 reg311,
                 reg310,
                 reg309,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 forvar298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 forvar293,
                 forvar292,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 forvar284,
                 reg283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 forvar278,
                 forvar277,
                 reg276,
                 reg275,
                 reg274,
                 reg273,
                 forvar272,
                 forvar271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 forvar264,
                 reg263,
                 reg262,
                 forvar261,
                 reg260,
                 forvar259,
                 reg258,
                 forvar257,
                 wire256,
                 wire255,
                 wire254,
                 wire252,
                 wire79,
                 wire78,
                 (1'h0)};
  assign wire78 = (+(^~(^wire77)));
  assign wire79 = (("ygCGL6rCICSL6Qk0HnQe" && wire78) ?
                      "6krB" : (($unsigned(wire78[(2'h2):(1'h0)]) ?
                          ({wire78} ?
                              (8'h9f) : {wire75}) : $unsigned($signed(wire76))) || wire75[(1'h1):(1'h0)]));
  module80 modinst253 (.clk(clk), .wire83(wire77), .wire82(wire78), .wire81(wire79), .y(wire252), .wire84(wire74));
  assign wire254 = (wire75 != (&wire76[(3'h4):(3'h4)]));
  assign wire255 = $unsigned(wire77[(3'h4):(3'h4)]);
  assign wire256 = $unsigned($unsigned((&($signed(wire77) ?
                       $signed(wire78) : {(8'ha4)}))));
  always
    @(posedge clk) begin
      for (forvar257 = (1'h0); (forvar257 < (1'h1)); forvar257 = (forvar257 + (1'h1)))
        begin
          reg258 <= ($signed(((wire78[(4'hb):(4'hb)] ?
                  $signed(wire76) : $unsigned((8'hb2))) ?
              (!wire74[(3'h6):(2'h3)]) : (^~(wire78 == wire74)))) ^ (-$unsigned((wire74[(3'h5):(3'h4)] & ((8'ha7) ?
              wire255 : wire256)))));
          for (forvar259 = (1'h0); (forvar259 < (2'h3)); forvar259 = (forvar259 + (1'h1)))
            begin
              reg260 = forvar257[(1'h1):(1'h0)];
            end
        end
      for (forvar261 = (1'h0); (forvar261 < (1'h0)); forvar261 = (forvar261 + (1'h1)))
        begin
          reg262 <= $unsigned((!$unsigned((+{wire255}))));
        end
      reg263 <= (-("qEouFW9l" > $unsigned(reg262)));
      for (forvar264 = (1'h0); (forvar264 < (1'h1)); forvar264 = (forvar264 + (1'h1)))
        begin
          reg265 <= $unsigned($unsigned($unsigned(wire75)));
          if ((!"xw9Xbvg"))
            begin
              reg266 <= (~&wire77[(2'h3):(1'h0)]);
            end
          else
            begin
              reg266 <= wire74[(3'h4):(3'h4)];
              reg267 = ((^{$unsigned($unsigned(forvar261)),
                  (~^((8'hab) < wire254))}) | ("dOSefyUv0aX" ?
                  (&forvar261[(1'h0):(1'h0)]) : $unsigned(($unsigned(forvar261) ?
                      (wire74 ? wire76 : reg260) : $signed((8'hbd))))));
              reg268 <= forvar264[(2'h3):(1'h1)];
            end
          if ({((reg267[(1'h0):(1'h0)] - "IYgGfA3bl3GMdMkrS3k") ?
                  "whmFpTG8eFDHt2bdo98t" : wire76)})
            begin
              reg269 <= (|(($signed((!wire252)) ?
                  $unsigned(forvar261[(2'h2):(2'h2)]) : reg262) | $signed($unsigned(reg260))));
              reg270 = {(8'hab)};
            end
          else
            begin
              reg269 = "bxP4QuAlMtDKc";
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar271 = (1'h0); (forvar271 < (1'h0)); forvar271 = (forvar271 + (1'h1)))
        begin
          for (forvar272 = (1'h0); (forvar272 < (1'h1)); forvar272 = (forvar272 + (1'h1)))
            begin
              reg273 <= {(reg268 ?
                      wire74[(3'h4):(2'h2)] : reg262[(4'ha):(3'h4)]),
                  $signed(forvar261)};
              reg274 <= $signed((^~($signed((8'h9f)) ?
                  $unsigned(reg263) : {(^~reg258)})));
              reg275 <= ($signed($signed({{forvar264, forvar272},
                  (+reg266)})) <<< (~&((((8'ha6) ?
                  reg263 : wire255) >> (reg268 ?
                  wire256 : wire78)) == $signed(reg262[(4'ha):(2'h2)]))));
            end
          reg276 <= wire75[(1'h1):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar277 = (1'h0); (forvar277 < (2'h3)); forvar277 = (forvar277 + (1'h1)))
        begin
          for (forvar278 = (1'h0); (forvar278 < (1'h0)); forvar278 = (forvar278 + (1'h1)))
            begin
              reg279 <= (!(8'ha9));
              reg280 <= $signed($unsigned($unsigned((wire79[(1'h0):(1'h0)] ?
                  (forvar272 ? (8'hac) : forvar278) : wire78))));
              reg281 <= (~&(~&{(!reg274)}));
              reg282 = ((8'h9d) ?
                  $unsigned((8'hb5)) : forvar257[(1'h0):(1'h0)]);
            end
          reg283 <= (|reg270[(3'h7):(3'h6)]);
          for (forvar284 = (1'h0); (forvar284 < (2'h3)); forvar284 = (forvar284 + (1'h1)))
            begin
              reg285 = ($signed($unsigned($signed(reg282[(3'h4):(1'h0)]))) ?
                  $unsigned(forvar284) : reg276[(4'h8):(2'h3)]);
              reg286 <= $signed($signed(({$signed(wire79)} ^~ {$unsigned(forvar278),
                  (reg275 > (8'h9d))})));
              reg287 = $unsigned((~(($signed(forvar277) <= (reg265 ^ (7'h43))) ?
                  {(^~forvar278), reg266} : (^~(reg285 ?
                      (8'hb4) : forvar259)))));
              reg288 <= wire75[(4'h9):(2'h2)];
              reg289 = $unsigned($unsigned($signed("pGVzY45I2p")));
            end
          reg290 <= (reg289 ?
              forvar277 : (forvar284 << (forvar272 ?
                  $signed($signed(reg279)) : (reg267[(1'h0):(1'h0)] <= (reg288 ?
                      (8'haa) : forvar257)))));
          reg291 = $unsigned($signed(reg262));
        end
      for (forvar292 = (1'h0); (forvar292 < (2'h3)); forvar292 = (forvar292 + (1'h1)))
        begin
          for (forvar293 = (1'h0); (forvar293 < (1'h1)); forvar293 = (forvar293 + (1'h1)))
            begin
              reg294 <= (reg289[(3'h4):(1'h1)] || ($unsigned(wire254) != (((^~wire78) <<< $unsigned(reg291)) ?
                  (~(reg258 ? reg260 : forvar272)) : {(~&wire78),
                      $signed(reg283)})));
              reg295 <= $signed((^~(+$unsigned($signed(reg276)))));
              reg296 = (7'h41);
              reg297 = (~&{forvar277});
            end
          for (forvar298 = (1'h0); (forvar298 < (3'h4)); forvar298 = (forvar298 + (1'h1)))
            begin
              reg299 <= $unsigned((($unsigned({forvar257, reg260}) ?
                      ((&(7'h42)) ?
                          $unsigned(reg297) : (wire255 | reg290)) : wire75) ?
                  (&$signed($unsigned((8'haf)))) : ($unsigned($signed(wire76)) ?
                      "DkFJWtf" : $unsigned((^reg273)))));
            end
          if ((-forvar277))
            begin
              reg300 <= (8'ha2);
              reg301 <= $signed($unsigned((({wire252,
                  forvar293} + $unsigned(reg296)) >>> "kGEDiy5hfSU2zzMq")));
              reg302 <= (wire74[(3'h7):(1'h0)] ?
                  $signed($signed(({reg265,
                      (7'h41)} >> (|forvar272)))) : reg269);
              reg303 <= reg301[(2'h3):(1'h0)];
              reg304 <= ((^~reg276) || reg299[(3'h7):(3'h6)]);
            end
          else
            begin
              reg300 <= ((reg282[(5'h11):(2'h2)] | $unsigned($signed($unsigned((8'hbe))))) ?
                  $signed($signed(($signed(forvar257) > (reg303 ?
                      reg287 : reg268)))) : $unsigned($signed(forvar271[(2'h3):(2'h3)])));
              reg301 <= $unsigned("205kw5rTh");
              reg302 <= forvar259;
            end
          if ($signed($signed((8'ha4))))
            begin
              reg305 <= wire76[(1'h0):(1'h0)];
              reg306 <= ({$signed(reg289)} << $unsigned($signed(((forvar298 ~^ forvar298) ^~ $unsigned(wire77)))));
              reg307 = $unsigned((~|$unsigned(reg295[(3'h4):(1'h1)])));
              reg308 = reg282;
              reg309 = (^(($unsigned({forvar272}) ~^ (&$unsigned(wire74))) && reg267));
            end
          else
            begin
              reg305 <= "kVm";
              reg306 <= ($unsigned(reg300[(4'hd):(3'h7)]) ?
                  $signed($unsigned((-(~forvar293)))) : ($unsigned($unsigned($signed(reg262))) + ((^forvar278[(1'h1):(1'h1)]) ?
                      {$unsigned(reg273), (reg294 ^ (8'h9d))} : ((wire252 ?
                              reg266 : (8'haf)) ?
                          reg301 : $unsigned(wire77)))));
            end
        end
      reg310 = $signed(forvar278);
    end
  always
    @(posedge clk) begin
      reg311 <= wire255[(3'h5):(3'h5)];
    end
  assign wire312 = (reg308 ? wire74[(3'h5):(1'h1)] : forvar272);
  module313 modinst435 (.wire316(forvar272), .y(wire434), .wire317(reg303), .clk(clk), .wire315(reg281), .wire314(reg270));
  always
    @(posedge clk) begin
      for (forvar436 = (1'h0); (forvar436 < (1'h0)); forvar436 = (forvar436 + (1'h1)))
        begin
          if ((wire76[(2'h2):(2'h2)] ?
              $unsigned((~^reg306[(3'h5):(3'h5)])) : {(forvar259[(2'h2):(2'h2)] ?
                      (|reg289[(4'h9):(3'h6)]) : {$unsigned((7'h44))})}))
            begin
              reg437 <= wire256;
            end
          else
            begin
              reg437 = ((^~"2KIa") ?
                  reg302 : ($signed($signed((8'hbc))) ?
                      wire76[(1'h0):(1'h0)] : reg279));
              reg438 <= $unsigned($signed({(8'hae), reg286[(1'h1):(1'h0)]}));
              reg439 = $signed((reg290[(5'h11):(4'hf)] || $signed("IqitkigV")));
            end
        end
      for (forvar440 = (1'h0); (forvar440 < (1'h0)); forvar440 = (forvar440 + (1'h1)))
        begin
          if ($signed($signed(((^~(~&reg288)) ?
              $unsigned(reg274[(2'h3):(1'h1)]) : $signed(reg299)))))
            begin
              reg441 = "JSGmhn";
              reg442 = {wire252[(5'h12):(3'h5)], $unsigned(reg297)};
              reg443 <= ((^wire76) ?
                  (|$unsigned((^{(8'hb9)}))) : $signed((((~(8'hba)) ?
                      $unsigned(reg266) : (8'hb5)) != $signed(reg283[(1'h1):(1'h1)]))));
            end
          else
            begin
              reg441 <= {(8'hb9)};
              reg442 = (^reg273[(4'ha):(2'h2)]);
              reg443 <= reg276[(3'h4):(1'h1)];
              reg444 = $unsigned(($signed($unsigned((reg301 ?
                  reg290 : reg443))) - ($signed($signed(reg260)) ^~ {(|reg296),
                  $signed(forvar278)})));
              reg445 = {(~({(reg263 - reg438)} >>> ((wire79 ?
                          forvar257 : reg279) ?
                      $unsigned(reg437) : reg269)))};
            end
          if ($unsigned({forvar298}))
            begin
              reg446 <= (~^(|(reg438 ~^ reg270)));
              reg447 = (~|$unsigned($unsigned($unsigned((reg441 - (8'ha5))))));
            end
          else
            begin
              reg446 <= (forvar440[(3'h6):(1'h1)] >= ($unsigned(reg310) ?
                  (reg305 ?
                      (&reg291) : (~$unsigned(reg308))) : ((|$unsigned(reg446)) ?
                      forvar271 : $signed((~|forvar271)))));
              reg447 = "hu5c37GIGle";
              reg448 = $signed({(reg300 && (+(reg267 <= (8'hbe)))),
                  $signed(forvar278)});
            end
          for (forvar449 = (1'h0); (forvar449 < (1'h1)); forvar449 = (forvar449 + (1'h1)))
            begin
              reg450 <= $signed(($signed(((-forvar436) ?
                      ((8'h9f) || wire256) : (~|reg446))) ?
                  {reg279,
                      reg305[(3'h6):(2'h3)]} : $signed($signed(reg263[(4'hd):(3'h5)]))));
            end
          if (($unsigned(wire79[(3'h5):(1'h1)]) == $signed((((reg276 ?
                  (8'hae) : wire76) & (wire74 ^ reg276)) ?
              ((-reg307) >>> wire75[(2'h3):(1'h1)]) : ((wire76 ?
                      (8'hb1) : reg280) ?
                  "" : $unsigned((8'ha1)))))))
            begin
              reg451 <= $unsigned(reg306);
              reg452 <= $unsigned(({reg301} >> {$unsigned($unsigned(forvar259))}));
            end
          else
            begin
              reg451 = ({($unsigned({reg295}) ?
                      "Snl7" : ($signed(reg302) ^ wire434))} <= (("1rtbvqhZSECkEw8KImR3" ?
                      ((-reg438) ?
                          forvar293 : reg439[(1'h1):(1'h1)]) : $unsigned(wire79[(2'h2):(2'h2)])) ?
                  (8'hb1) : (~^((~|reg437) >> ((8'hba) ?
                      forvar259 : reg258)))));
              reg452 <= (8'had);
              reg453 <= $signed($unsigned(wire254[(3'h4):(1'h0)]));
            end
        end
      reg454 <= $signed($signed(((~|forvar440[(1'h1):(1'h0)]) + (~|$signed(reg263)))));
    end
  always
    @(posedge clk) begin
      reg455 <= (reg441 ?
          "ep0KRr" : $unsigned((reg438[(4'h8):(2'h2)] ?
              (8'ha1) : (~&$unsigned(reg270)))));
      reg456 = $unsigned(("NakNCwDJbruyJE" & reg309[(4'h8):(3'h4)]));
      for (forvar457 = (1'h0); (forvar457 < (2'h2)); forvar457 = (forvar457 + (1'h1)))
        begin
          reg458 <= reg304[(3'h4):(1'h0)];
          for (forvar459 = (1'h0); (forvar459 < (2'h3)); forvar459 = (forvar459 + (1'h1)))
            begin
              reg460 <= ((!({(reg301 <= reg446)} ?
                      (~&(!forvar264)) : $signed((-(8'hbf))))) ?
                  $signed(reg262) : (reg263 ?
                      (|(reg438[(3'h4):(2'h3)] ?
                          wire312[(4'h8):(2'h2)] : reg456[(1'h1):(1'h0)])) : $unsigned(reg265[(3'h6):(3'h6)])));
              reg461 = (+(^(((|reg273) ?
                  (reg279 | reg275) : $unsigned(forvar259)) ~^ $signed(reg452))));
              reg462 = ((^{($unsigned((8'ha7)) >> (~|wire77))}) ?
                  reg268[(2'h2):(1'h1)] : wire255[(4'hc):(2'h2)]);
              reg463 <= $unsigned((-$signed($signed((8'haa)))));
              reg464 <= $signed(reg454[(3'h7):(1'h1)]);
            end
          reg465 <= $signed((!(({reg262, forvar271} ?
                  ((8'hbd) < reg446) : $unsigned(forvar272)) ?
              (~&{(8'had)}) : reg455[(2'h3):(2'h2)])));
          reg466 <= $signed((($unsigned(wire76[(1'h1):(1'h0)]) <<< (~&$unsigned(forvar440))) | (8'ha4)));
          reg467 <= (((reg306[(4'hf):(4'hf)] && (^(+reg267))) ?
                  $signed($unsigned($unsigned(reg437))) : reg282) ?
              reg307 : $signed(reg301));
        end
      reg468 <= reg296[(1'h1):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg469 <= $signed(reg263[(3'h7):(3'h7)]);
      for (forvar470 = (1'h0); (forvar470 < (1'h0)); forvar470 = (forvar470 + (1'h1)))
        begin
          if (reg466[(2'h2):(1'h1)])
            begin
              reg471 = reg453[(4'h9):(4'h9)];
              reg472 <= reg294;
            end
          else
            begin
              reg471 = reg307[(3'h5):(3'h4)];
              reg472 <= (!{((^(~&reg444)) != (8'hb2))});
              reg473 = {reg285[(2'h2):(2'h2)], reg303};
              reg474 = ((($signed(reg300) ?
                      $unsigned($signed(reg283)) : reg448) ^~ "byRX2QCTHhDyYET") ?
                  (~^reg466[(1'h1):(1'h0)]) : reg467[(2'h3):(1'h0)]);
              reg475 = $unsigned((($unsigned((reg268 ?
                      reg286 : (8'ha8))) == forvar293) ?
                  reg263[(4'hb):(3'h4)] : {(~^(forvar261 == reg447))}));
            end
          for (forvar476 = (1'h0); (forvar476 < (1'h1)); forvar476 = (forvar476 + (1'h1)))
            begin
              reg477 = reg307;
              reg478 <= reg311;
            end
          reg479 <= ($signed(wire256[(4'hd):(1'h1)]) ^ (+reg441));
          if ((($unsigned($signed((&reg463))) ?
                  reg295[(4'h9):(2'h3)] : (reg444[(4'hb):(4'ha)] == (((8'ha1) <= forvar470) && (forvar449 ?
                      reg276 : reg305)))) ?
              (&reg475) : reg454[(2'h3):(2'h3)]))
            begin
              reg480 = $unsigned($unsigned(reg269[(2'h2):(2'h2)]));
              reg481 <= ({($signed((8'had)) <= (|(~|reg450)))} ?
                  (|(reg308[(2'h3):(1'h0)] * reg475[(5'h12):(4'h8)])) : (((~&reg282[(3'h5):(1'h1)]) ?
                          (reg288[(1'h1):(1'h1)] >>> reg473[(4'hc):(4'hb)]) : ("bFVuluG0dQMlHxTa9ND9" & reg297[(1'h0):(1'h0)])) ?
                      reg475 : $signed((~|(forvar277 - reg468)))));
            end
          else
            begin
              reg480 = (!(~|(+$signed(wire312))));
              reg481 <= ((reg471 ?
                  $signed($signed($signed(reg296))) : {$unsigned($signed(reg269))}) >> $unsigned(reg306));
              reg482 = (((reg451 <<< $signed(reg291[(2'h2):(2'h2)])) >= $unsigned($signed(reg307))) ?
                  (forvar298[(1'h0):(1'h0)] >= reg471) : reg442);
              reg483 <= (~((^$signed(reg285[(2'h3):(2'h2)])) >> (^~(8'had))));
            end
        end
    end
  assign wire484 = (8'hba);
  assign wire485 = ($unsigned($signed(($signed(wire78) ?
                           $unsigned(forvar278) : $unsigned(reg280)))) ?
                       ((forvar440 ?
                               reg291[(3'h4):(2'h2)] : ((reg479 | reg441) & $signed(reg477))) ?
                           (reg453[(3'h5):(1'h1)] - reg304[(2'h3):(2'h2)]) : reg468[(1'h0):(1'h0)]) : reg437);
  assign wire486 = $unsigned((($unsigned(reg445) ?
                       $signed((~|wire434)) : ((8'hae) < reg280[(1'h0):(1'h0)])) >= forvar436[(2'h2):(1'h0)]));
  assign wire487 = reg309;
  assign wire488 = reg460;
  assign wire489 = $unsigned(reg285);
  assign wire490 = (reg280 <= wire488);
  assign wire491 = (~&(wire490 ? (!reg469) : wire255[(1'h0):(1'h0)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module313
#( parameter param432 = (~&(!(~^(((8'ha6) >= (8'ha8)) ? ((8'h9c) ? (8'h9e) : (7'h43)) : ((8'hab) ? (7'h42) : (8'ha8))))))
, parameter param433 = param432 )
(y, clk, wire317, wire316, wire315, wire314);
  output wire [(32'h540):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire317;
  input wire signed [(5'h12):(1'h0)] wire316;
  input wire signed [(2'h3):(1'h0)] wire315;
  input wire signed [(4'he):(1'h0)] wire314;
  wire signed [(4'ha):(1'h0)] wire431;
  reg signed [(3'h6):(1'h0)] reg430 = (1'h0);
  reg [(4'hd):(1'h0)] reg429 = (1'h0);
  reg [(5'h13):(1'h0)] forvar428 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg427 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg426 = (1'h0);
  reg [(5'h13):(1'h0)] reg425 = (1'h0);
  reg [(3'h6):(1'h0)] forvar424 = (1'h0);
  reg [(3'h6):(1'h0)] reg423 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg422 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg421 = (1'h0);
  reg [(4'ha):(1'h0)] reg420 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg419 = (1'h0);
  reg [(5'h13):(1'h0)] reg418 = (1'h0);
  reg [(5'h15):(1'h0)] reg417 = (1'h0);
  reg [(3'h7):(1'h0)] reg416 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg415 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar414 = (1'h0);
  reg [(5'h10):(1'h0)] forvar413 = (1'h0);
  reg [(3'h5):(1'h0)] reg412 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg401 = (1'h0);
  reg [(3'h6):(1'h0)] forvar398 = (1'h0);
  reg [(5'h11):(1'h0)] reg397 = (1'h0);
  reg [(4'hb):(1'h0)] reg395 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg411 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg410 = (1'h0);
  reg [(5'h13):(1'h0)] reg409 = (1'h0);
  reg [(4'he):(1'h0)] reg408 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg407 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar406 = (1'h0);
  reg [(5'h15):(1'h0)] reg405 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg404 = (1'h0);
  reg [(4'hb):(1'h0)] reg403 = (1'h0);
  reg [(3'h6):(1'h0)] reg402 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar401 = (1'h0);
  reg [(4'h8):(1'h0)] reg400 = (1'h0);
  reg [(3'h6):(1'h0)] reg399 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg398 = (1'h0);
  reg [(5'h13):(1'h0)] forvar397 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg396 = (1'h0);
  reg [(2'h3):(1'h0)] forvar395 = (1'h0);
  reg signed [(4'he):(1'h0)] reg394 = (1'h0);
  reg [(3'h4):(1'h0)] reg393 = (1'h0);
  wire [(3'h5):(1'h0)] wire392;
  wire signed [(4'hf):(1'h0)] wire391;
  wire signed [(5'h14):(1'h0)] wire390;
  wire signed [(3'h6):(1'h0)] wire389;
  wire [(4'ha):(1'h0)] wire388;
  reg signed [(5'h12):(1'h0)] reg387 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg386 = (1'h0);
  reg [(5'h13):(1'h0)] forvar385 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg384 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg383 = (1'h0);
  wire [(2'h3):(1'h0)] wire382;
  reg [(3'h7):(1'h0)] reg381 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg380 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg379 = (1'h0);
  reg [(5'h11):(1'h0)] reg378 = (1'h0);
  reg [(4'he):(1'h0)] reg377 = (1'h0);
  reg [(4'hb):(1'h0)] forvar376 = (1'h0);
  reg [(4'h8):(1'h0)] forvar375 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg374 = (1'h0);
  reg [(4'h9):(1'h0)] reg373 = (1'h0);
  reg [(4'h9):(1'h0)] reg372 = (1'h0);
  reg signed [(4'he):(1'h0)] reg371 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar370 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar369 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg368 = (1'h0);
  reg [(4'h8):(1'h0)] forvar367 = (1'h0);
  wire [(4'h8):(1'h0)] wire366;
  wire [(4'hf):(1'h0)] wire365;
  wire signed [(5'h14):(1'h0)] wire364;
  wire signed [(3'h6):(1'h0)] wire363;
  wire [(4'hf):(1'h0)] wire362;
  wire signed [(5'h12):(1'h0)] wire361;
  reg [(3'h6):(1'h0)] reg360 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg359 = (1'h0);
  wire [(4'hc):(1'h0)] wire358;
  wire signed [(4'hd):(1'h0)] wire357;
  reg signed [(3'h4):(1'h0)] reg356 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg355 = (1'h0);
  reg signed [(4'he):(1'h0)] reg354 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg353 = (1'h0);
  reg [(4'hf):(1'h0)] reg352 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg351 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg350 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar349 = (1'h0);
  reg signed [(4'he):(1'h0)] reg348 = (1'h0);
  reg [(3'h4):(1'h0)] reg347 = (1'h0);
  reg [(2'h2):(1'h0)] reg346 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg345 = (1'h0);
  reg [(4'hf):(1'h0)] reg344 = (1'h0);
  reg [(2'h3):(1'h0)] forvar343 = (1'h0);
  reg [(2'h2):(1'h0)] forvar342 = (1'h0);
  reg [(2'h3):(1'h0)] forvar325 = (1'h0);
  reg [(4'h8):(1'h0)] reg324 = (1'h0);
  reg [(4'hc):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg340 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar339 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg338 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg337 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg336 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg335 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg334 = (1'h0);
  reg [(3'h4):(1'h0)] reg333 = (1'h0);
  reg [(5'h12):(1'h0)] reg332 = (1'h0);
  reg [(5'h10):(1'h0)] reg331 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar330 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg329 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg328 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg327 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg326 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg325 = (1'h0);
  reg [(3'h6):(1'h0)] forvar324 = (1'h0);
  reg [(5'h12):(1'h0)] reg323 = (1'h0);
  reg [(4'h9):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg321 = (1'h0);
  reg [(4'he):(1'h0)] reg320 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg319 = (1'h0);
  reg [(4'h9):(1'h0)] forvar318 = (1'h0);
  assign y = {wire431,
                 reg430,
                 reg429,
                 forvar428,
                 reg427,
                 reg426,
                 reg425,
                 forvar424,
                 reg423,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 forvar414,
                 forvar413,
                 reg412,
                 reg401,
                 forvar398,
                 reg397,
                 reg395,
                 reg411,
                 reg410,
                 reg409,
                 reg408,
                 reg407,
                 forvar406,
                 reg405,
                 reg404,
                 reg403,
                 reg402,
                 forvar401,
                 reg400,
                 reg399,
                 reg398,
                 forvar397,
                 reg396,
                 forvar395,
                 reg394,
                 reg393,
                 wire392,
                 wire391,
                 wire390,
                 wire389,
                 wire388,
                 reg387,
                 reg386,
                 forvar385,
                 reg384,
                 reg383,
                 wire382,
                 reg381,
                 reg380,
                 reg379,
                 reg378,
                 reg377,
                 forvar376,
                 forvar375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 forvar370,
                 forvar369,
                 reg368,
                 forvar367,
                 wire366,
                 wire365,
                 wire364,
                 wire363,
                 wire362,
                 wire361,
                 reg360,
                 reg359,
                 wire358,
                 wire357,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 reg351,
                 reg350,
                 forvar349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg344,
                 forvar343,
                 forvar342,
                 forvar325,
                 reg324,
                 reg341,
                 reg340,
                 forvar339,
                 reg338,
                 reg337,
                 reg336,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg331,
                 forvar330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 forvar324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 forvar318,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (($signed($signed($unsigned($unsigned(wire314)))) >= ((~|{$signed(wire317),
          $unsigned(wire314)}) > wire315)))
        begin
          for (forvar318 = (1'h0); (forvar318 < (3'h4)); forvar318 = (forvar318 + (1'h1)))
            begin
              reg319 <= ((&$unsigned({(!wire316), $unsigned(wire314)})) ?
                  wire315 : (+wire314[(1'h0):(1'h0)]));
              reg320 <= (8'had);
              reg321 <= $signed($signed({$signed((!wire314))}));
              reg322 <= (|wire314[(3'h7):(1'h1)]);
              reg323 <= $signed(((((~&wire315) | wire315[(1'h1):(1'h1)]) <= {(reg320 ?
                          reg319 : wire316),
                      reg320}) ?
                  "dOyM9JV3H64g7KZG" : {{(^~reg321), wire315}}));
            end
          for (forvar324 = (1'h0); (forvar324 < (1'h1)); forvar324 = (forvar324 + (1'h1)))
            begin
              reg325 <= ($signed(((&"7NvQZMuS0PK0kFK2Bp") ?
                      ((~wire316) ?
                          $signed(forvar324) : reg321) : (~&reg323[(4'hb):(1'h0)]))) ?
                  ((({wire314} ?
                          reg322[(1'h1):(1'h1)] : reg320[(3'h6):(1'h1)]) ?
                      "zfWq5w8habErfCp9Oht" : (8'hae)) >> (~&($unsigned(wire315) ?
                      (forvar324 + reg323) : $signed(wire316)))) : ((&(~|$unsigned((7'h42)))) | $signed(($signed((8'ha4)) ?
                      (^forvar318) : (&wire315)))));
              reg326 = $unsigned(($unsigned($unsigned((wire317 ?
                  reg321 : wire317))) ~^ reg322[(3'h4):(2'h2)]));
              reg327 = (~reg325);
              reg328 <= $unsigned(reg320[(3'h6):(3'h5)]);
              reg329 <= ({$unsigned((reg328[(4'he):(1'h0)] & {reg323})),
                  {$signed(forvar318[(3'h5):(3'h4)])}} * "hhNifl8holfOMsX");
            end
          for (forvar330 = (1'h0); (forvar330 < (2'h3)); forvar330 = (forvar330 + (1'h1)))
            begin
              reg331 <= ({reg325[(3'h6):(2'h3)]} ?
                  {(wire317[(3'h6):(2'h2)] ?
                          $signed($signed((7'h42))) : (forvar318[(2'h3):(2'h2)] ?
                              {wire314, wire314} : $unsigned(wire314))),
                      $unsigned($signed(((8'ha3) & reg322)))} : ((8'ha5) ?
                      (((-(8'hbc)) ?
                          reg328[(4'h9):(4'h8)] : (reg327 >= wire314)) == ($signed((8'ha2)) * $unsigned((8'haf)))) : (wire315 - (8'ha3))));
              reg332 = (!{((wire317[(4'ha):(3'h7)] < $signed(wire314)) < $unsigned((~&forvar330)))});
              reg333 <= ((reg331[(4'hd):(3'h5)] ^ ({$signed((8'hb3)),
                      (reg331 ^ forvar324)} > $unsigned(reg323[(4'hf):(4'ha)]))) ?
                  (8'ha2) : forvar318[(1'h1):(1'h0)]);
              reg334 <= forvar324;
            end
          if ("iI")
            begin
              reg335 = ($signed($unsigned({reg328[(4'he):(4'hb)]})) ?
                  $signed((forvar318 & (~|$signed(reg327)))) : reg327[(4'ha):(4'h9)]);
              reg336 = (8'hab);
              reg337 <= ($unsigned(((~&$signed(reg331)) ?
                      $unsigned((~|reg332)) : wire315[(1'h0):(1'h0)])) ?
                  ((((+wire317) <<< (reg326 ? reg333 : forvar318)) ?
                      reg325 : ($unsigned(reg321) ?
                          (reg329 ?
                              reg319 : reg333) : reg336)) <= reg327[(1'h0):(1'h0)]) : (reg320[(4'hd):(3'h5)] || {($signed((7'h41)) & $signed(reg336)),
                      {wire316, wire314[(4'ha):(1'h1)]}}));
            end
          else
            begin
              reg335 <= reg331;
              reg336 = (~^$signed(reg334));
              reg337 <= (reg323[(5'h11):(5'h11)] || reg323[(2'h3):(1'h0)]);
              reg338 <= $unsigned($unsigned(forvar324));
            end
          for (forvar339 = (1'h0); (forvar339 < (1'h1)); forvar339 = (forvar339 + (1'h1)))
            begin
              reg340 <= ("PWQR7ruehw6afWH" ?
                  ((-$signed(reg331[(3'h7):(3'h7)])) && ((8'had) && forvar324[(3'h4):(1'h0)])) : reg333);
              reg341 <= reg334;
            end
        end
      else
        begin
          for (forvar318 = (1'h0); (forvar318 < (2'h3)); forvar318 = (forvar318 + (1'h1)))
            begin
              reg319 <= (reg322[(3'h6):(2'h2)] * reg327);
              reg320 = (($signed(wire315[(2'h2):(1'h0)]) ?
                      reg333 : reg335[(2'h3):(2'h2)]) ?
                  (~|(8'hbb)) : reg336[(4'hc):(4'hc)]);
              reg321 <= reg332[(4'h8):(3'h5)];
              reg322 = reg325[(2'h3):(1'h1)];
              reg323 <= $signed(reg335);
            end
          reg324 <= $unsigned($unsigned(("HiHIP3klzav3OOw4o" ?
              reg336[(3'h6):(2'h3)] : (|{(8'hb8), (8'hbc)}))));
          for (forvar325 = (1'h0); (forvar325 < (1'h1)); forvar325 = (forvar325 + (1'h1)))
            begin
              reg326 = (~(^~(($signed(reg326) <<< (-reg333)) ?
                  wire316 : (7'h43))));
            end
        end
      for (forvar342 = (1'h0); (forvar342 < (1'h1)); forvar342 = (forvar342 + (1'h1)))
        begin
          for (forvar343 = (1'h0); (forvar343 < (2'h3)); forvar343 = (forvar343 + (1'h1)))
            begin
              reg344 <= $signed(forvar318[(3'h5):(2'h3)]);
              reg345 = (reg324[(1'h1):(1'h1)] ?
                  ((-{$unsigned(forvar324), reg337[(2'h3):(2'h3)]}) ?
                      reg321 : ($unsigned((7'h41)) ?
                          ({reg340, reg323} && (forvar339 ?
                              reg328 : reg338)) : $signed($unsigned((8'h9f))))) : forvar339);
              reg346 = reg345[(4'hc):(4'ha)];
              reg347 = $signed(forvar318[(2'h2):(2'h2)]);
              reg348 <= reg325[(4'h9):(4'h9)];
            end
          for (forvar349 = (1'h0); (forvar349 < (1'h1)); forvar349 = (forvar349 + (1'h1)))
            begin
              reg350 <= reg321;
            end
          reg351 <= $unsigned(("ciGK3xSwJVQsc6a" ?
              $signed((|(forvar349 ^ (8'h9d)))) : {"iuT6A8",
                  $unsigned((+reg337))}));
          if ($unsigned(forvar325))
            begin
              reg352 = (+(forvar324 ? $signed(reg333[(2'h3):(1'h0)]) : reg332));
              reg353 <= $signed(reg350);
              reg354 <= $signed(reg351[(1'h0):(1'h0)]);
              reg355 <= (8'hac);
              reg356 <= reg326[(2'h2):(1'h0)];
            end
          else
            begin
              reg352 = reg332[(4'h9):(1'h0)];
            end
        end
    end
  assign wire357 = ((($signed($unsigned(reg321)) << (((8'ha1) ?
                           reg341 : reg334) ?
                       (reg324 ? reg344 : forvar325) : (reg323 ?
                           (8'ha8) : forvar330))) ~^ (~reg334[(2'h2):(1'h1)])) >= (^~$signed((~|{(8'ha4),
                       forvar339}))));
  assign wire358 = (-{$unsigned(reg335)});
  always
    @(posedge clk) begin
      reg359 <= (|$signed(forvar318[(4'h9):(3'h4)]));
      reg360 = (-$signed(((~|(forvar349 * wire357)) <= reg345)));
    end
  assign wire361 = (~$unsigned(forvar339[(2'h3):(2'h3)]));
  assign wire362 = {wire317, reg345[(1'h1):(1'h0)]};
  assign wire363 = $unsigned((wire314 | (forvar349[(3'h4):(2'h2)] ?
                       reg354[(4'h8):(3'h5)] : reg346[(1'h1):(1'h1)])));
  assign wire364 = wire316[(4'hc):(1'h1)];
  assign wire365 = (((~"3MWNcwF2") ?
                           "YSsgA" : $unsigned($unsigned($unsigned(reg335)))) ?
                       ($unsigned(("4RSHCqmKeNEHs" <= (!reg340))) - (^~reg336[(4'h8):(3'h4)])) : $signed(((+"7aURtC6JM7obMcynSWH") ?
                           (reg348[(1'h1):(1'h1)] ?
                               (~&reg356) : ((8'ha9) ?
                                   (8'ha0) : reg346)) : $unsigned(((8'hbf) <= forvar324)))));
  assign wire366 = $unsigned($signed({wire361, reg354}));
  always
    @(posedge clk) begin
      for (forvar367 = (1'h0); (forvar367 < (2'h3)); forvar367 = (forvar367 + (1'h1)))
        begin
          if ($signed(((~{(^reg344)}) || $signed("QYYnRZQZZ"))))
            begin
              reg368 = ((^(((+(8'ha3)) ? wire366 : $signed((8'hb7))) ?
                      {$signed(reg360),
                          reg335[(3'h4):(1'h0)]} : (forvar330[(4'h9):(3'h5)] >= wire366))) ?
                  (+((reg332[(1'h0):(1'h0)] ?
                          {reg331, forvar342} : "ZZCmIfSosg9u2I") ?
                      $unsigned(((7'h40) || reg335)) : $unsigned($unsigned(reg324)))) : ((|wire315) ?
                      $unsigned((~$signed(reg350))) : reg335[(2'h2):(1'h0)]));
            end
          else
            begin
              reg368 = (^~{(reg329 >>> $signed($unsigned(reg344))), forvar324});
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar369 = (1'h0); (forvar369 < (2'h3)); forvar369 = (forvar369 + (1'h1)))
        begin
          for (forvar370 = (1'h0); (forvar370 < (2'h3)); forvar370 = (forvar370 + (1'h1)))
            begin
              reg371 = $signed((-(forvar325[(2'h3):(2'h3)] ?
                  $unsigned((8'h9d)) : reg332)));
              reg372 = ((~(&(reg344 || {wire314, wire364}))) ?
                  $signed(reg320[(1'h1):(1'h1)]) : (8'hbf));
              reg373 = (reg353 ?
                  (($unsigned((reg336 == wire362)) >>> $unsigned(reg338)) || reg344) : "vFgrR9i");
              reg374 <= "PLdmk";
            end
        end
      for (forvar375 = (1'h0); (forvar375 < (2'h2)); forvar375 = (forvar375 + (1'h1)))
        begin
          for (forvar376 = (1'h0); (forvar376 < (3'h4)); forvar376 = (forvar376 + (1'h1)))
            begin
              reg377 <= reg371;
              reg378 <= wire317[(4'h9):(3'h7)];
            end
          if ((((~|((~&reg336) ?
              {wire314} : {(8'ha1)})) <= ($unsigned($signed((8'haf))) * $signed(reg378))) == ((reg335[(1'h1):(1'h0)] >>> reg377[(4'h8):(2'h2)]) << (reg331[(4'hc):(3'h7)] && wire363))))
            begin
              reg379 <= {$unsigned((!forvar370[(1'h1):(1'h0)])),
                  ($unsigned({((8'h9c) <<< wire316)}) ?
                      reg378[(5'h11):(4'h8)] : ($unsigned(reg337) ?
                          reg337[(4'h9):(4'h9)] : (wire357[(4'ha):(2'h2)] | $signed(reg320))))};
              reg380 = $unsigned((|{forvar349[(1'h0):(1'h0)],
                  (^~reg323[(3'h5):(1'h0)])}));
            end
          else
            begin
              reg379 <= $signed((^$signed((reg331 ?
                  ((8'hb2) >> reg327) : $unsigned(reg352)))));
              reg380 = (reg371 ?
                  $unsigned(((8'ha0) ^ ((^~reg335) ?
                      ((8'hbd) ~^ (7'h41)) : $signed((8'hb4))))) : $signed((+(~&(wire365 ?
                      (8'h9f) : forvar369)))));
            end
          reg381 <= reg377;
        end
    end
  assign wire382 = ($unsigned((~|$signed(reg359[(3'h6):(1'h1)]))) == ($signed($signed((-(8'hae)))) ?
                       {(~reg373[(3'h4):(2'h2)]),
                           ((forvar370 ? wire364 : reg338) ?
                               reg335[(3'h4):(1'h0)] : $signed(reg353))} : ({(reg346 >> reg341)} ?
                           $unsigned($signed(reg335)) : {(^reg346),
                               (reg380 ? forvar367 : reg374)})));
  always
    @(posedge clk) begin
      reg383 <= reg338;
      reg384 <= $unsigned(wire358);
      for (forvar385 = (1'h0); (forvar385 < (1'h0)); forvar385 = (forvar385 + (1'h1)))
        begin
          reg386 <= forvar330;
          reg387 = $unsigned((8'hb0));
        end
    end
  assign wire388 = $signed({$signed(({reg323} ?
                           (reg344 == reg324) : ((7'h41) ? wire363 : (8'hab)))),
                       $unsigned(((reg380 >>> forvar367) >>> (~&reg346)))});
  assign wire389 = (+{((|(wire365 | (8'hae))) + (^(reg341 || wire366)))});
  assign wire390 = {((~&$signed($signed(reg329))) | ($signed((~&reg344)) ?
                           $unsigned(reg338) : (reg360[(3'h6):(2'h2)] << (reg321 ?
                               wire314 : reg378))))};
  assign wire391 = reg379;
  assign wire392 = reg341;
  always
    @(posedge clk) begin
      reg393 <= $unsigned(reg321);
      if ($signed($signed($signed((+(reg374 ? reg380 : reg377))))))
        begin
          reg394 = ((+"C0") ? wire314 : reg319[(1'h0):(1'h0)]);
          for (forvar395 = (1'h0); (forvar395 < (3'h4)); forvar395 = (forvar395 + (1'h1)))
            begin
              reg396 <= "2lKfUF0";
            end
          for (forvar397 = (1'h0); (forvar397 < (1'h1)); forvar397 = (forvar397 + (1'h1)))
            begin
              reg398 <= reg326;
              reg399 <= (("3lQRa321uT1Q" ?
                  reg352 : "nf6gKCVTkrS1bb3vX") < wire365[(3'h4):(1'h0)]);
              reg400 = (&(~&{((&forvar367) <= reg327[(3'h7):(3'h4)])}));
            end
          for (forvar401 = (1'h0); (forvar401 < (1'h1)); forvar401 = (forvar401 + (1'h1)))
            begin
              reg402 <= ((!(-$signed(wire390))) ?
                  reg324[(3'h7):(1'h0)] : $unsigned(wire364[(4'h9):(2'h3)]));
              reg403 <= $signed(((reg378[(2'h2):(1'h0)] ?
                  (^~(reg384 ?
                      reg386 : (8'hbf))) : $unsigned((-(7'h41)))) && ""));
              reg404 = $signed(("sthnTamLwwg" ?
                  forvar397 : (~$unsigned(reg331[(2'h2):(1'h1)]))));
              reg405 = (8'h9d);
            end
          for (forvar406 = (1'h0); (forvar406 < (2'h3)); forvar406 = (forvar406 + (1'h1)))
            begin
              reg407 = (($signed($signed(wire389)) + reg394) ?
                  $unsigned(forvar324[(1'h0):(1'h0)]) : {($signed((-reg378)) ?
                          ($signed(forvar375) > $unsigned(wire358)) : wire314[(3'h6):(3'h5)])});
              reg408 <= (8'h9c);
              reg409 <= reg344;
              reg410 = (^(~|(($unsigned((8'hae)) ?
                  (-reg320) : (reg384 == reg332)) == $signed($unsigned(wire365)))));
              reg411 <= ((~|{(reg319 ? (+(8'hb8)) : $unsigned(wire364))}) ?
                  $signed(reg393) : (^$unsigned(({forvar375} ?
                      "" : $signed(reg331)))));
            end
        end
      else
        begin
          reg394 <= reg332[(5'h10):(1'h1)];
          if (($unsigned(reg329[(3'h6):(3'h6)]) ?
              ((^~$unsigned($unsigned(forvar406))) ?
                  $unsigned($signed($signed(forvar397))) : wire363[(2'h2):(1'h0)]) : $unsigned(($signed(reg398) ?
                  ($unsigned(reg394) <<< (~^reg384)) : (+(reg384 ?
                      reg368 : wire314))))))
            begin
              reg395 <= $unsigned($signed(reg410));
              reg396 <= $unsigned(($unsigned($unsigned($signed((8'hb2)))) ^~ reg387[(1'h1):(1'h1)]));
            end
          else
            begin
              reg395 = wire391;
              reg396 = (^($unsigned((~|reg333)) ?
                  reg338[(4'hd):(3'h5)] : {((8'hb4) ? (~^reg333) : {reg340}),
                      ((8'haa) ?
                          (~^reg400) : (forvar370 ? wire361 : reg359))}));
              reg397 <= reg387[(1'h0):(1'h0)];
            end
          for (forvar398 = (1'h0); (forvar398 < (1'h1)); forvar398 = (forvar398 + (1'h1)))
            begin
              reg399 <= $signed((&((&reg340) ?
                  {(8'hb1)} : $signed(wire314[(2'h2):(1'h0)]))));
              reg400 <= reg395[(4'hb):(1'h0)];
              reg401 <= (+(reg394[(4'he):(4'hd)] ?
                  ($signed(wire391) ^ ($signed(reg334) <<< (reg410 * (8'hbe)))) : forvar339));
              reg402 <= (|($signed(wire314) ?
                  reg332[(3'h5):(1'h1)] : ($signed("") <= ((reg322 - reg334) ?
                      $unsigned(forvar406) : $signed(reg380)))));
            end
          reg403 = $unsigned((~|$signed(((&reg325) ?
              {(8'hba)} : $unsigned(forvar330)))));
          reg404 = $unsigned((reg331 ?
              ({{(8'hac), (7'h44)}} && reg386) : wire316));
        end
      reg412 <= ((|(((!reg368) & wire314[(2'h3):(1'h0)]) < ((forvar342 ?
              reg374 : reg324) != wire358[(3'h4):(1'h0)]))) ?
          (~"Q1W") : $unsigned((reg380[(2'h2):(1'h1)] - ((7'h41) > (reg352 | forvar376)))));
      for (forvar413 = (1'h0); (forvar413 < (2'h2)); forvar413 = (forvar413 + (1'h1)))
        begin
          for (forvar414 = (1'h0); (forvar414 < (2'h2)); forvar414 = (forvar414 + (1'h1)))
            begin
              reg415 = (wire358 ?
                  $signed(((~^$unsigned(reg380)) ?
                      {$unsigned(forvar330)} : "PnoU0SwyrKqC")) : reg324[(3'h7):(1'h0)]);
              reg416 = {(reg381[(3'h6):(2'h2)] ?
                      reg404 : $signed((wire366[(2'h2):(1'h0)] ?
                          $signed(reg393) : (reg384 != wire362))))};
              reg417 <= (($unsigned((forvar339[(3'h6):(1'h1)] * $unsigned(reg338))) ^ ((reg403[(4'h9):(4'h8)] ?
                      {reg345} : ((8'ha9) ? reg351 : wire366)) ?
                  reg372 : reg393[(3'h4):(1'h0)])) <<< $unsigned($unsigned(((-wire389) ?
                  $unsigned(reg398) : $unsigned(reg404)))));
              reg418 <= $unsigned("hW0ZbHXtdG4g");
              reg419 <= {wire315[(2'h3):(1'h1)], (!forvar406[(3'h6):(1'h1)])};
            end
          reg420 = (~&($unsigned($signed($signed(forvar367))) * reg403));
          if ($unsigned((&(($signed(reg401) + reg328[(4'hb):(2'h3)]) & {(^~reg395),
              (~wire362)}))))
            begin
              reg421 <= ({reg396[(3'h6):(3'h6)],
                      (+((reg403 ? reg331 : reg360) > (!wire316)))} ?
                  ((8'ha3) ?
                      $unsigned(($signed((8'hba)) || (!reg386))) : ((~wire364) <<< reg374)) : (^~((((8'hb0) ?
                          reg335 : forvar376) + (~|forvar375)) ?
                      (&(^~reg394)) : $signed(forvar406))));
              reg422 = $unsigned((~|forvar325));
            end
          else
            begin
              reg421 <= {(~^(|reg359))};
              reg422 <= $unsigned((forvar318[(3'h5):(3'h4)] ^ wire382[(2'h3):(1'h0)]));
              reg423 <= wire390;
            end
          for (forvar424 = (1'h0); (forvar424 < (2'h3)); forvar424 = (forvar424 + (1'h1)))
            begin
              reg425 <= (reg321[(4'hd):(4'ha)] <<< (((~forvar370) ?
                  (+reg412[(2'h3):(1'h0)]) : $unsigned(reg351)) >>> $unsigned((~&((8'hbb) ?
                  (8'h9f) : reg359)))));
              reg426 <= ($signed($signed(forvar406[(1'h1):(1'h0)])) & $signed(wire364));
              reg427 <= (8'hb7);
            end
          for (forvar428 = (1'h0); (forvar428 < (3'h4)); forvar428 = (forvar428 + (1'h1)))
            begin
              reg429 <= reg355;
            end
        end
      reg430 = {(8'hb3)};
    end
  assign wire431 = $unsigned(reg355);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module80
#( parameter param251 = ((!(!(((8'ha4) ^ (7'h44)) || ((8'hb3) ? (8'ha0) : (7'h42))))) ? ((|((~|(8'h9d)) + (~|(7'h40)))) ? (+(((8'hae) ? (8'ha0) : (8'ha0)) ? ((8'h9c) ? (8'ha2) : (8'hbc)) : ((8'ha0) ? (8'hb8) : (8'had)))) : (8'hbb)) : (((((8'hbd) ? (8'hb3) : (8'h9f)) ? ((8'h9d) ? (8'hb3) : (8'hb0)) : (^~(8'hac))) ? {((8'h9e) ? (8'ha4) : (8'hae)), (~^(8'haf))} : (((8'ha2) ~^ (8'ha5)) ? ((8'hac) >>> (8'ha7)) : (~(8'ha8)))) ? (({(8'hb1)} + (~&(7'h42))) ? ((!(8'ha2)) || (+(8'hb8))) : (((7'h44) && (8'ha0)) && ((8'hb3) ? (8'h9f) : (8'hb8)))) : ((~^(|(8'hbc))) ? (&{(8'hbe)}) : {((7'h42) ? (8'ha1) : (8'haa)), ((8'ha9) >= (8'hb4))}))) )
(y, clk, wire84, wire83, wire82, wire81);
  output wire [(32'h792):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire84;
  input wire [(4'h8):(1'h0)] wire83;
  input wire [(4'he):(1'h0)] wire82;
  input wire [(4'hc):(1'h0)] wire81;
  wire signed [(4'hd):(1'h0)] wire250;
  reg [(5'h11):(1'h0)] reg249 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg248 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg247 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg246 = (1'h0);
  reg [(4'ha):(1'h0)] reg245 = (1'h0);
  reg [(5'h12):(1'h0)] forvar244 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg243 = (1'h0);
  reg [(5'h10):(1'h0)] reg242 = (1'h0);
  reg [(5'h12):(1'h0)] reg241 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg240 = (1'h0);
  reg [(2'h2):(1'h0)] reg239 = (1'h0);
  reg [(5'h13):(1'h0)] forvar238 = (1'h0);
  reg [(4'h9):(1'h0)] reg237 = (1'h0);
  reg [(4'ha):(1'h0)] reg236 = (1'h0);
  reg [(4'hd):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar233 = (1'h0);
  reg [(2'h3):(1'h0)] forvar232 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire231;
  wire signed [(4'hb):(1'h0)] wire230;
  wire signed [(5'h10):(1'h0)] wire229;
  wire signed [(4'h9):(1'h0)] wire228;
  wire [(4'h8):(1'h0)] wire227;
  reg signed [(3'h5):(1'h0)] reg226 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg225 = (1'h0);
  reg [(4'hd):(1'h0)] reg224 = (1'h0);
  reg [(4'h8):(1'h0)] reg223 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg222 = (1'h0);
  reg [(3'h6):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg220 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg219 = (1'h0);
  reg [(5'h13):(1'h0)] reg218 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg212 = (1'h0);
  reg [(2'h3):(1'h0)] reg217 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg216 = (1'h0);
  reg [(5'h14):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg214 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg213 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar212 = (1'h0);
  reg [(4'hd):(1'h0)] reg211 = (1'h0);
  reg [(5'h13):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar209 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg208 = (1'h0);
  reg [(5'h15):(1'h0)] reg207 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg195 = (1'h0);
  reg [(5'h12):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg205 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg204 = (1'h0);
  reg [(3'h4):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg202 = (1'h0);
  reg [(4'hc):(1'h0)] forvar201 = (1'h0);
  reg [(3'h5):(1'h0)] reg200 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg199 = (1'h0);
  reg [(3'h6):(1'h0)] reg198 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg197 = (1'h0);
  reg [(4'ha):(1'h0)] reg196 = (1'h0);
  reg [(4'ha):(1'h0)] forvar195 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg194 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg193 = (1'h0);
  reg [(3'h6):(1'h0)] reg192 = (1'h0);
  reg [(4'he):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg190 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg189 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg188 = (1'h0);
  reg [(3'h5):(1'h0)] reg187 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar186 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg185 = (1'h0);
  reg [(5'h14):(1'h0)] reg184 = (1'h0);
  reg [(3'h7):(1'h0)] reg183 = (1'h0);
  reg [(4'hb):(1'h0)] reg182 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar181 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg181 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg180 = (1'h0);
  reg [(4'hd):(1'h0)] reg179 = (1'h0);
  reg [(2'h2):(1'h0)] reg178 = (1'h0);
  reg [(4'hb):(1'h0)] forvar177 = (1'h0);
  reg [(5'h13):(1'h0)] reg176 = (1'h0);
  reg [(3'h5):(1'h0)] reg175 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg174 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg173 = (1'h0);
  reg [(4'he):(1'h0)] reg172 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar171 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar170 = (1'h0);
  reg [(2'h3):(1'h0)] reg169 = (1'h0);
  wire [(3'h6):(1'h0)] wire168;
  reg signed [(5'h11):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg166 = (1'h0);
  reg [(4'h9):(1'h0)] reg165 = (1'h0);
  reg [(5'h14):(1'h0)] forvar164 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg163 = (1'h0);
  reg [(3'h7):(1'h0)] reg162 = (1'h0);
  reg [(3'h5):(1'h0)] reg161 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg160 = (1'h0);
  reg [(3'h5):(1'h0)] forvar159 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg158 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg157 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg156 = (1'h0);
  reg [(3'h4):(1'h0)] reg155 = (1'h0);
  reg [(3'h7):(1'h0)] forvar154 = (1'h0);
  reg [(4'he):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg152 = (1'h0);
  reg [(4'he):(1'h0)] reg151 = (1'h0);
  reg [(5'h10):(1'h0)] reg150 = (1'h0);
  reg [(4'h9):(1'h0)] reg149 = (1'h0);
  reg [(4'h8):(1'h0)] forvar148 = (1'h0);
  reg [(5'h11):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg146 = (1'h0);
  reg [(3'h6):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg144 = (1'h0);
  reg [(4'h9):(1'h0)] reg143 = (1'h0);
  reg [(3'h7):(1'h0)] reg142 = (1'h0);
  reg [(3'h7):(1'h0)] reg141 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg140 = (1'h0);
  reg [(5'h15):(1'h0)] reg139 = (1'h0);
  reg [(4'hc):(1'h0)] reg138 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar137 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar136 = (1'h0);
  reg [(4'ha):(1'h0)] reg135 = (1'h0);
  reg [(5'h11):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg133 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar132 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar131 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg117 = (1'h0);
  reg [(5'h10):(1'h0)] reg130 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg129 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg127 = (1'h0);
  reg [(4'h8):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg125 = (1'h0);
  reg [(2'h2):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar123 = (1'h0);
  reg [(5'h10):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg121 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg120 = (1'h0);
  reg [(5'h11):(1'h0)] reg119 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg118 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar117 = (1'h0);
  reg [(5'h12):(1'h0)] reg116 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg115 = (1'h0);
  reg [(4'he):(1'h0)] reg114 = (1'h0);
  reg [(5'h14):(1'h0)] reg113 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar112 = (1'h0);
  reg [(3'h5):(1'h0)] reg111 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg106 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg103 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg110 = (1'h0);
  reg [(4'hc):(1'h0)] reg109 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg108 = (1'h0);
  reg [(4'ha):(1'h0)] reg107 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar106 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg105 = (1'h0);
  reg [(2'h3):(1'h0)] reg104 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar103 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg102 = (1'h0);
  reg [(2'h2):(1'h0)] reg101 = (1'h0);
  reg [(5'h11):(1'h0)] forvar100 = (1'h0);
  reg [(5'h14):(1'h0)] reg99 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg98 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg97 = (1'h0);
  reg [(4'hd):(1'h0)] reg96 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg95 = (1'h0);
  reg [(3'h6):(1'h0)] reg94 = (1'h0);
  reg [(5'h14):(1'h0)] reg93 = (1'h0);
  reg [(4'he):(1'h0)] reg92 = (1'h0);
  reg [(4'h9):(1'h0)] reg91 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg90 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg89 = (1'h0);
  reg [(5'h11):(1'h0)] forvar88 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg87 = (1'h0);
  reg [(4'hd):(1'h0)] forvar86 = (1'h0);
  wire [(4'ha):(1'h0)] wire85;
  assign y = {wire250,
                 reg249,
                 reg248,
                 reg247,
                 reg246,
                 reg245,
                 forvar244,
                 reg243,
                 reg242,
                 reg241,
                 reg240,
                 reg239,
                 forvar238,
                 reg237,
                 reg236,
                 reg235,
                 reg234,
                 forvar233,
                 forvar232,
                 wire231,
                 wire230,
                 wire229,
                 wire228,
                 wire227,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 reg212,
                 reg217,
                 reg216,
                 reg215,
                 reg214,
                 reg213,
                 forvar212,
                 reg211,
                 reg210,
                 forvar209,
                 reg208,
                 reg207,
                 reg195,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 forvar201,
                 reg200,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 forvar195,
                 reg194,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 forvar186,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 forvar181,
                 reg181,
                 reg180,
                 reg179,
                 reg178,
                 forvar177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg172,
                 forvar171,
                 forvar170,
                 reg169,
                 wire168,
                 reg167,
                 reg166,
                 reg165,
                 forvar164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 forvar159,
                 reg158,
                 reg157,
                 reg156,
                 reg155,
                 forvar154,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 forvar148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 forvar137,
                 forvar136,
                 reg135,
                 reg134,
                 reg133,
                 forvar132,
                 forvar131,
                 reg117,
                 reg130,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 forvar123,
                 reg122,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 forvar117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 forvar112,
                 reg111,
                 reg106,
                 reg103,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 forvar106,
                 reg105,
                 reg104,
                 forvar103,
                 reg102,
                 reg101,
                 forvar100,
                 reg99,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 forvar88,
                 reg87,
                 forvar86,
                 wire85,
                 (1'h0)};
  assign wire85 = (~{($unsigned((wire82 ? wire84 : wire81)) ?
                          ((wire84 || wire81) ?
                              $unsigned((8'hba)) : wire81) : (~|(wire84 <= wire81)))});
  always
    @(posedge clk) begin
      for (forvar86 = (1'h0); (forvar86 < (2'h3)); forvar86 = (forvar86 + (1'h1)))
        begin
          reg87 <= (~wire85[(4'ha):(2'h3)]);
          for (forvar88 = (1'h0); (forvar88 < (1'h1)); forvar88 = (forvar88 + (1'h1)))
            begin
              reg89 = wire83;
              reg90 <= (~&wire84);
              reg91 <= wire82;
              reg92 <= wire83;
            end
          reg93 <= {(~^((forvar86 >>> $signed((8'hbe))) ?
                  (reg87[(5'h15):(5'h10)] <= wire83) : forvar86)),
              (~&reg90[(2'h2):(1'h1)])};
          if ($signed(((~^wire84) ?
              ({(wire82 ?
                      wire82 : (8'h9c))} >>> ((|forvar88) ~^ forvar86[(3'h5):(1'h0)])) : ((reg93[(4'ha):(1'h1)] ?
                      $signed(wire83) : (reg92 ^ reg90)) ?
                  $unsigned((~&wire84)) : $unsigned(wire81[(4'hb):(3'h6)])))))
            begin
              reg94 <= $signed($unsigned(wire82[(4'h9):(1'h1)]));
              reg95 <= reg91;
              reg96 = $unsigned(reg94[(1'h0):(1'h0)]);
              reg97 = (~^wire85);
            end
          else
            begin
              reg94 <= (&$signed(((^~$signed(wire83)) > wire84)));
              reg95 <= $signed($unsigned(reg93));
              reg96 <= (reg96[(2'h2):(2'h2)] ?
                  $unsigned((8'h9c)) : (wire84[(4'h8):(3'h5)] >>> ($unsigned((reg87 <<< reg94)) >>> ((8'hbd) ?
                      (forvar88 | wire83) : (~|reg94)))));
            end
          reg98 <= $unsigned((7'h42));
        end
      reg99 <= (reg90 ?
          {"ZR5txNn26ugqmqwyQiL",
              wire82[(1'h0):(1'h0)]} : reg91[(1'h1):(1'h0)]);
      for (forvar100 = (1'h0); (forvar100 < (2'h3)); forvar100 = (forvar100 + (1'h1)))
        begin
          reg101 <= "pVfghcFr3wcKTxY";
          reg102 <= forvar86[(4'hc):(4'hb)];
        end
    end
  always
    @(posedge clk) begin
      if ({(!$signed($signed((forvar88 * reg89))))})
        begin
          for (forvar103 = (1'h0); (forvar103 < (3'h4)); forvar103 = (forvar103 + (1'h1)))
            begin
              reg104 <= (reg99 ? reg89 : "n9");
              reg105 <= reg91;
            end
          for (forvar106 = (1'h0); (forvar106 < (2'h3)); forvar106 = (forvar106 + (1'h1)))
            begin
              reg107 = "brnGRvKc";
              reg108 = {{(reg87[(5'h14):(5'h11)] != $unsigned((reg95 + reg105))),
                      {($unsigned((8'ha0)) ? wire84[(2'h3):(2'h3)] : (8'ha9)),
                          reg98}},
                  reg87[(1'h1):(1'h1)]};
            end
          reg109 = $signed(((forvar106[(3'h6):(3'h6)] ?
              reg90[(3'h6):(3'h5)] : (|(~|(8'h9e)))) ~^ ($signed($signed(reg97)) ?
              forvar103 : $unsigned((8'hb1)))));
          reg110 = (|(8'hbd));
        end
      else
        begin
          reg103 = {wire81[(4'ha):(3'h6)], reg101};
          reg104 <= (^~$unsigned(($signed({(7'h42),
              forvar86}) >> {$signed(reg104)})));
          reg105 = reg91[(1'h0):(1'h0)];
          reg106 <= ({"CxYQOnuAbqlq2ZEt",
              ($unsigned($signed(reg97)) < $signed({reg99}))} <= ($signed({(~&reg96)}) ?
              (+("NiVl4" > ((8'ha1) ?
                  wire84 : reg108))) : $unsigned(reg87[(5'h11):(4'he)])));
        end
      reg111 = ((~&(!$unsigned({(8'hb9)}))) >> (!reg93[(4'hc):(4'hb)]));
      for (forvar112 = (1'h0); (forvar112 < (2'h2)); forvar112 = (forvar112 + (1'h1)))
        begin
          if (reg98[(4'h9):(3'h5)])
            begin
              reg113 = $signed($signed($signed($signed((reg107 >>> forvar103)))));
            end
          else
            begin
              reg113 <= (reg103[(5'h13):(3'h6)] ?
                  ({$signed($signed(reg101))} ^ (forvar106 ?
                      reg113[(4'h9):(3'h7)] : ($unsigned(forvar106) ^~ (wire85 ?
                          forvar106 : reg87)))) : ($unsigned(("5QJBNmJFyEFMC4O0KMNy" ?
                      (reg90 ?
                          (8'ha2) : reg92) : reg102[(3'h7):(3'h5)])) ~^ reg103));
              reg114 <= (8'hac);
              reg115 = {reg96,
                  ((~&(wire81 + $signed(reg107))) ?
                      (reg107[(2'h2):(2'h2)] ?
                          (8'hbc) : $unsigned((~|reg94))) : (~^forvar103[(4'h9):(4'h8)]))};
              reg116 <= reg94;
            end
        end
    end
  always
    @(posedge clk) begin
      if ((($signed(reg98) ?
          reg98[(1'h0):(1'h0)] : ($unsigned($signed(reg97)) || $signed({(8'hb1),
              reg101}))) < ($signed(reg92) ?
          reg95[(4'h9):(4'h8)] : (+$unsigned($signed(reg99))))))
        begin
          for (forvar117 = (1'h0); (forvar117 < (2'h3)); forvar117 = (forvar117 + (1'h1)))
            begin
              reg118 <= reg105[(3'h5):(2'h2)];
              reg119 <= {reg90, $signed($signed(reg98))};
              reg120 = (&($unsigned($signed((reg107 ?
                  reg96 : wire81))) | ({reg91} ?
                  forvar112[(1'h1):(1'h0)] : (+{forvar103}))));
              reg121 <= (reg89[(1'h1):(1'h1)] ?
                  {$signed(forvar117)} : $signed($unsigned(forvar100[(4'hf):(3'h7)])));
              reg122 = (^reg104);
            end
          for (forvar123 = (1'h0); (forvar123 < (2'h2)); forvar123 = (forvar123 + (1'h1)))
            begin
              reg124 <= (~(^(~|(8'h9c))));
              reg125 <= reg101;
              reg126 <= (((((wire85 ? reg121 : wire84) - {forvar100, reg87}) ?
                          (forvar123 >= $unsigned(reg94)) : (~&reg125)) ?
                      forvar86[(4'hc):(2'h3)] : reg96[(4'ha):(2'h2)]) ?
                  {forvar112[(1'h0):(1'h0)],
                      (forvar123[(2'h3):(2'h3)] ?
                          {(|reg107),
                              (8'ha3)} : $unsigned(forvar88[(4'hf):(2'h3)]))} : ((!$signed(reg98)) ?
                      "GhMoqN1knWFh4Zuwe" : (reg91 ?
                          reg120 : $signed(forvar103))));
              reg127 = (reg96 ?
                  ((reg97[(2'h3):(2'h3)] >>> (+$signed(reg109))) >= $signed(wire85[(1'h0):(1'h0)])) : reg96[(4'hb):(1'h0)]);
            end
          reg128 <= ($signed($unsigned(reg119[(2'h3):(2'h2)])) ^ reg110);
          reg129 <= $signed((reg107[(4'h8):(3'h6)] ?
              $unsigned({$unsigned(reg92),
                  (reg89 ?
                      reg107 : reg126)}) : $unsigned(wire84[(3'h7):(3'h7)])));
          reg130 <= $unsigned(((^((wire83 ?
                  reg121 : wire82) ^ (reg109 - reg98))) ?
              $unsigned((((8'hb8) ? reg101 : reg110) ?
                  (reg116 ? reg125 : reg93) : {(8'ha3),
                      reg122})) : $signed(((reg128 > reg89) & ((8'ha7) ?
                  forvar112 : forvar117)))));
        end
      else
        begin
          reg117 <= (8'h9f);
        end
      for (forvar131 = (1'h0); (forvar131 < (2'h3)); forvar131 = (forvar131 + (1'h1)))
        begin
          for (forvar132 = (1'h0); (forvar132 < (2'h2)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 <= $signed((forvar100 ?
                  $unsigned(reg129[(3'h6):(3'h6)]) : $signed(reg120[(3'h4):(2'h2)])));
              reg134 = $unsigned(((($signed(forvar132) ?
                      reg120 : (forvar86 ^~ reg102)) && (~^$signed(reg91))) ?
                  ($unsigned($signed(reg102)) ^ (~^$unsigned(reg93))) : $signed({(~wire83),
                      reg124})));
              reg135 = "";
            end
        end
      for (forvar136 = (1'h0); (forvar136 < (2'h2)); forvar136 = (forvar136 + (1'h1)))
        begin
          for (forvar137 = (1'h0); (forvar137 < (1'h0)); forvar137 = (forvar137 + (1'h1)))
            begin
              reg138 <= (((|$signed((reg109 >>> reg91))) ?
                  $unsigned(forvar88) : (reg90[(3'h4):(3'h4)] >> reg129)) << reg133);
              reg139 = ({reg108[(3'h6):(1'h0)],
                      $signed((^~(reg89 ? reg118 : reg128)))} ?
                  reg116 : forvar117[(3'h4):(2'h2)]);
              reg140 = (reg134 ? (8'hb3) : $signed(reg126[(2'h3):(2'h3)]));
              reg141 = {(8'hb9)};
              reg142 <= $signed(reg92[(3'h5):(1'h0)]);
            end
          if ($signed((reg90[(3'h4):(1'h1)] >= (reg133 | ((&reg135) ^~ {reg130})))))
            begin
              reg143 = (8'hb0);
              reg144 = (reg135 ?
                  (~^$signed(forvar112[(2'h2):(1'h0)])) : (^~reg119));
              reg145 = reg124[(2'h2):(2'h2)];
              reg146 <= $unsigned({$signed(reg133),
                  ("z1UIWWq68gm" >> forvar112[(2'h3):(1'h0)])});
            end
          else
            begin
              reg143 <= ((!(~^reg120)) ?
                  {((reg102 <<< (reg90 ? reg145 : (8'haf))) || ((wire85 ?
                          reg124 : reg119) ^~ reg134))} : $signed($unsigned((reg113[(5'h14):(3'h6)] ?
                      ((7'h40) ? forvar100 : reg92) : ((8'ha6) ?
                          (8'hb1) : reg111)))));
              reg144 <= $signed(((~^{(&reg90)}) || {$unsigned((reg91 ?
                      reg117 : reg91)),
                  $signed((reg120 >> forvar86))}));
              reg145 <= ($signed("") - {$unsigned(reg140),
                  ((reg95 ? (reg110 * reg110) : $unsigned((8'hbe))) ?
                      $unsigned($unsigned(reg97)) : reg115)});
              reg146 <= $unsigned(($unsigned(({reg127, forvar112} >= reg143)) ?
                  (wire83[(4'h8):(1'h1)] ?
                      $unsigned((8'hb6)) : $signed(reg114[(3'h7):(3'h7)])) : $unsigned(reg103[(4'h9):(3'h4)])));
              reg147 <= (reg109 & (($signed({reg128, reg104}) ?
                  (~(forvar131 ?
                      reg104 : reg93)) : $signed((reg142 == (8'hbe)))) && (-($unsigned(reg101) ?
                  $signed(reg104) : {reg105}))));
            end
          for (forvar148 = (1'h0); (forvar148 < (2'h2)); forvar148 = (forvar148 + (1'h1)))
            begin
              reg149 <= (8'hae);
              reg150 = (reg125 << (~|$unsigned((~^reg143[(3'h6):(1'h1)]))));
              reg151 = $signed(($signed(wire81[(4'h9):(4'h9)]) ?
                  (8'hac) : $signed($signed(reg91[(2'h2):(1'h1)]))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg152 = ((8'hab) << $unsigned(((^~(reg94 ? forvar103 : reg120)) ?
          reg99 : ((reg113 <= (8'hab)) ?
              (reg122 ? (8'hb8) : forvar137) : (forvar137 ? reg97 : reg99)))));
      reg153 <= (reg149[(3'h6):(3'h5)] ?
          reg103[(1'h0):(1'h0)] : forvar131[(3'h4):(2'h2)]);
      for (forvar154 = (1'h0); (forvar154 < (3'h4)); forvar154 = (forvar154 + (1'h1)))
        begin
          reg155 = reg128[(1'h0):(1'h0)];
          reg156 <= {$signed((reg93[(5'h11):(1'h0)] ?
                  reg106[(3'h7):(3'h7)] : reg133))};
          reg157 <= $unsigned(("cllGol2Olok" ?
              wire84 : $unsigned(((reg106 && reg98) || reg117[(4'h8):(2'h2)]))));
        end
      reg158 = (wire82[(4'ha):(3'h4)] | $unsigned((($unsigned(reg134) ?
          $unsigned((8'hbe)) : reg113) <<< {{(8'hbb), reg99},
          ((7'h44) != reg87)})));
      for (forvar159 = (1'h0); (forvar159 < (1'h0)); forvar159 = (forvar159 + (1'h1)))
        begin
          reg160 <= $unsigned("ybz49bm0BqmLhpKqY");
          reg161 <= reg150;
          reg162 = reg160[(2'h2):(2'h2)];
          reg163 <= (^(reg130 << reg125[(5'h11):(2'h2)]));
          for (forvar164 = (1'h0); (forvar164 < (1'h0)); forvar164 = (forvar164 + (1'h1)))
            begin
              reg165 <= (^reg97[(3'h4):(3'h4)]);
              reg166 = {(($unsigned(reg156[(1'h1):(1'h0)]) < reg108[(1'h1):(1'h0)]) ?
                      forvar132 : ({(reg151 ? reg151 : reg110)} ?
                          {$unsigned(reg103)} : ((reg156 << reg113) ?
                              (reg157 * reg147) : (~&reg128)))),
                  (reg99 + (!$signed($signed(reg143))))};
              reg167 <= ($unsigned((reg90[(1'h1):(1'h0)] - {$signed(reg142),
                      $unsigned(reg163)})) ?
                  $unsigned($unsigned($unsigned(reg94[(3'h5):(1'h1)]))) : forvar136[(3'h5):(2'h3)]);
            end
        end
    end
  assign wire168 = reg153[(4'h9):(1'h1)];
  always
    @(posedge clk) begin
      reg169 = wire81;
      for (forvar170 = (1'h0); (forvar170 < (1'h0)); forvar170 = (forvar170 + (1'h1)))
        begin
          for (forvar171 = (1'h0); (forvar171 < (1'h0)); forvar171 = (forvar171 + (1'h1)))
            begin
              reg172 = $signed((8'hbe));
              reg173 = {$unsigned(wire81)};
              reg174 = reg169[(1'h1):(1'h0)];
              reg175 = (-forvar148);
            end
        end
      reg176 = $signed(reg139[(3'h5):(1'h1)]);
      if ($unsigned(($unsigned(reg107[(3'h4):(1'h1)]) ?
          reg172[(3'h7):(1'h0)] : forvar112[(2'h2):(2'h2)])))
        begin
          for (forvar177 = (1'h0); (forvar177 < (2'h2)); forvar177 = (forvar177 + (1'h1)))
            begin
              reg178 <= reg108;
              reg179 <= $signed(reg178);
              reg180 <= (|((((~|(8'hb7)) ?
                      $signed(reg91) : reg161[(3'h4):(3'h4)]) >>> (^((7'h40) == (7'h41)))) ?
                  reg113[(4'hb):(3'h6)] : reg165[(3'h4):(1'h0)]));
            end
          reg181 <= $unsigned(({$signed((&forvar170)),
              reg105} || ($signed($unsigned(reg118)) || (forvar86[(4'hc):(3'h6)] ?
              {reg146} : ((8'hac) ? forvar112 : (8'hbf))))));
        end
      else
        begin
          for (forvar177 = (1'h0); (forvar177 < (3'h4)); forvar177 = (forvar177 + (1'h1)))
            begin
              reg178 <= reg165;
            end
          reg179 = $signed((8'h9e));
          reg180 <= ($unsigned((~{reg146[(4'ha):(4'h9)]})) ?
              (!(!$unsigned((reg95 >>> reg174)))) : reg174);
          for (forvar181 = (1'h0); (forvar181 < (2'h2)); forvar181 = (forvar181 + (1'h1)))
            begin
              reg182 = {$unsigned((((~^wire85) ?
                          (|(8'hb9)) : (reg158 + (8'hb7))) ?
                      $signed((reg114 ?
                          forvar177 : reg89)) : (forvar177[(4'h8):(1'h0)] ?
                          $unsigned(reg160) : (forvar132 <= reg90)))),
                  ("u2qbo" * reg106[(1'h1):(1'h1)])};
              reg183 <= {(-(!$signed((reg179 ? forvar154 : reg182)))),
                  $signed($unsigned((reg133[(4'h8):(1'h1)] ?
                      (!(8'hb3)) : (&reg91))))};
              reg184 = (|$signed(reg155));
              reg185 <= reg90[(1'h1):(1'h0)];
            end
          for (forvar186 = (1'h0); (forvar186 < (2'h2)); forvar186 = (forvar186 + (1'h1)))
            begin
              reg187 <= $signed($signed({reg122[(4'hf):(3'h7)],
                  ((|reg145) || (8'h9f))}));
              reg188 = ((+$unsigned("NyRnJwCdlwk")) ?
                  {(+($unsigned((8'hbf)) != (wire83 >>> forvar123)))} : {reg117});
              reg189 <= $unsigned(reg96[(4'hd):(4'h8)]);
            end
        end
      if ($unsigned((-{{$signed(reg143), ((8'h9c) == forvar159)},
          $signed($signed(reg141))})))
        begin
          if ($signed($signed((-reg116))))
            begin
              reg190 <= {$signed($signed($unsigned((8'hbd)))),
                  reg105[(1'h1):(1'h1)]};
            end
          else
            begin
              reg190 <= ((~^(reg102 >= {{(8'haa)},
                  (reg146 ? forvar112 : reg189)})) >> reg149[(4'h9):(3'h4)]);
              reg191 = reg89[(1'h1):(1'h0)];
              reg192 <= reg145;
              reg193 = ($signed(forvar123[(4'h8):(2'h2)]) ~^ (("6yR333UpH4fEn3MmAWE4" && {{forvar112,
                          (8'hb8)}}) ?
                  ((((8'hb2) ? wire83 : wire82) ?
                          (reg111 ? reg152 : reg162) : (~reg121)) ?
                      $signed((reg122 ?
                          reg169 : reg130)) : (^~reg102)) : (8'hb3)));
              reg194 = $signed(($unsigned((^(~reg142))) ?
                  $unsigned(reg92) : $unsigned(reg193[(1'h0):(1'h0)])));
            end
          for (forvar195 = (1'h0); (forvar195 < (1'h1)); forvar195 = (forvar195 + (1'h1)))
            begin
              reg196 <= (+wire83[(1'h1):(1'h0)]);
              reg197 = reg190;
              reg198 = $signed((~&(|forvar100)));
              reg199 <= "Xoh1YrXEzoxeBEhl";
            end
          reg200 <= ((&reg183) ? reg89[(1'h1):(1'h1)] : forvar86);
          for (forvar201 = (1'h0); (forvar201 < (2'h3)); forvar201 = (forvar201 + (1'h1)))
            begin
              reg202 <= $unsigned((forvar164 == ($signed((-reg121)) ?
                  ($signed(forvar132) ?
                      reg129 : $unsigned(reg155)) : ((forvar103 < reg160) ?
                      {forvar177} : $unsigned(forvar117)))));
              reg203 <= ((~&(reg149 ^~ forvar106)) && (-(($unsigned(reg167) <= (&forvar148)) ?
                  $unsigned("HOpo3Y") : (8'haa))));
              reg204 <= forvar137[(4'hd):(1'h0)];
              reg205 = $signed($signed(($signed(reg193) ?
                  reg197 : reg176[(5'h13):(5'h13)])));
              reg206 <= (((~&((|reg129) >> (~|wire168))) ?
                  ($unsigned((~reg97)) + "R1GU") : $unsigned(reg180)) != reg188);
            end
        end
      else
        begin
          if ($signed($unsigned(reg175[(3'h4):(1'h1)])))
            begin
              reg190 <= $signed($signed((({wire82, forvar186} > {reg157,
                      reg94}) ?
                  (reg141[(1'h0):(1'h0)] || reg174[(2'h2):(1'h0)]) : $signed($signed(forvar106)))));
              reg191 <= reg118[(2'h3):(1'h1)];
              reg192 <= {(~&(!{$unsigned(forvar186)}))};
              reg193 <= reg188[(3'h6):(2'h3)];
              reg194 <= $signed($unsigned(("QMeCCKSTqHgsaG" << (~(reg126 ?
                  (8'hb9) : reg141)))));
            end
          else
            begin
              reg190 = ($signed((&((reg95 ?
                  reg197 : reg152) << reg105))) - $unsigned((wire168[(3'h4):(2'h2)] <= (^~((8'ha7) ?
                  reg134 : reg142)))));
              reg191 = forvar117[(4'h9):(3'h7)];
              reg192 = reg101[(1'h0):(1'h0)];
            end
          reg195 = reg203;
        end
    end
  always
    @(posedge clk) begin
      reg207 = ($unsigned(reg110) >> (~|(~^$unsigned($unsigned(forvar177)))));
      reg208 <= (^((^{$unsigned(reg141)}) ^ (((reg144 ?
              reg165 : reg199) <<< $unsigned(reg206)) ?
          {reg133[(4'ha):(3'h5)], (8'hb2)} : $unsigned((~wire81)))));
      for (forvar209 = (1'h0); (forvar209 < (2'h2)); forvar209 = (forvar209 + (1'h1)))
        begin
          reg210 = ({$signed((~^(-reg101)))} >= ({{reg105[(1'h0):(1'h0)],
                      (reg156 ? reg121 : forvar159)},
                  (^~wire168[(2'h3):(2'h3)])} ?
              (reg139 && reg202[(4'h8):(3'h5)]) : $signed((~^reg199))));
        end
      reg211 <= ((reg204[(5'h11):(4'he)] ?
          {$unsigned({forvar132})} : reg114) * (8'hb3));
    end
  always
    @(posedge clk) begin
      if ($signed($signed($unsigned(((~^(8'hbf)) ?
          (8'ha4) : ((8'hb7) < reg97))))))
        begin
          for (forvar212 = (1'h0); (forvar212 < (2'h3)); forvar212 = (forvar212 + (1'h1)))
            begin
              reg213 <= (~^forvar195);
              reg214 <= "GmQp";
              reg215 = ($signed({$unsigned(reg95)}) ?
                  $signed(reg101) : $signed(reg162[(1'h1):(1'h1)]));
              reg216 = (-($signed({$unsigned((8'ha2)),
                  reg173[(2'h3):(1'h1)]}) >>> ((reg195 ?
                  forvar100[(5'h10):(4'h9)] : (reg206 ?
                      reg151 : reg120)) << wire84[(3'h6):(3'h6)])));
            end
          reg217 = (~&{$unsigned($unsigned(reg214))});
        end
      else
        begin
          reg212 <= (^~($signed((reg216 > reg125[(4'hf):(1'h1)])) ^~ (8'hae)));
          if ($unsigned($signed(reg139[(1'h1):(1'h0)])))
            begin
              reg213 <= ($signed($unsigned(reg199[(4'h9):(4'h9)])) >> ((-reg146[(5'h10):(4'h9)]) ~^ (~(+reg93))));
              reg214 <= (reg90[(3'h4):(2'h2)] ? reg143 : reg90);
              reg215 = {reg188[(3'h5):(2'h3)]};
              reg216 <= reg105[(4'hb):(1'h0)];
            end
          else
            begin
              reg213 <= $signed(reg161[(1'h0):(1'h0)]);
              reg214 <= ("tVvJ3dvQvbrH7PEsBp" + reg145[(1'h0):(1'h0)]);
              reg215 <= (8'ha8);
            end
          reg217 <= forvar88;
          reg218 = (7'h44);
          if ((-$unsigned((~^$unsigned(reg94)))))
            begin
              reg219 = reg133;
              reg220 = (reg141 != $signed(reg202));
              reg221 = reg141[(3'h6):(3'h5)];
              reg222 <= (((({reg130} ? (|forvar181) : {reg206, reg144}) ?
                          reg175[(2'h3):(2'h3)] : ((~|reg162) - reg125)) ?
                      reg204 : "Qaf4qJt5kSuOffRhSP") ?
                  reg99 : $signed((|$signed({reg175}))));
              reg223 <= ({$unsigned(($unsigned(reg121) + reg138[(4'h9):(1'h1)])),
                  reg193} < (8'hb2));
            end
          else
            begin
              reg219 <= reg213[(5'h12):(5'h11)];
              reg220 <= {reg221[(1'h1):(1'h1)], $signed(reg188[(4'h8):(3'h7)])};
            end
        end
    end
  always
    @(posedge clk) begin
      reg224 <= $unsigned($signed((-reg139)));
      reg225 = $signed(reg93[(5'h14):(5'h12)]);
      reg226 = reg163[(2'h3):(2'h3)];
    end
  assign wire227 = (reg93 ?
                       $signed(($signed($unsigned(reg158)) ?
                           reg111[(3'h4):(3'h4)] : (reg129 <<< (reg203 ?
                               wire85 : wire85)))) : reg110[(1'h1):(1'h0)]);
  assign wire228 = reg183;
  assign wire229 = $signed((~&(reg158 && reg116)));
  assign wire230 = reg182[(4'ha):(1'h1)];
  assign wire231 = {reg125};
  always
    @(posedge clk) begin
      for (forvar232 = (1'h0); (forvar232 < (2'h2)); forvar232 = (forvar232 + (1'h1)))
        begin
          for (forvar233 = (1'h0); (forvar233 < (2'h3)); forvar233 = (forvar233 + (1'h1)))
            begin
              reg234 = (^~"5RFRLNfGsbiYUCx8nA");
              reg235 <= ($unsigned(wire229[(3'h7):(3'h7)]) | (reg181[(3'h4):(2'h3)] ?
                  ((8'ha4) * ((8'hb8) ?
                      $signed((8'h9d)) : forvar112[(1'h1):(1'h0)])) : (reg198[(3'h5):(3'h4)] * "zBq9KOZb1VYWC2pxCOwz")));
              reg236 <= reg149[(1'h1):(1'h0)];
              reg237 = ((&($signed(reg101[(1'h1):(1'h1)]) && (((8'hb0) + wire229) ?
                  (reg146 <<< forvar181) : (reg150 && (8'hb2))))) || forvar117);
            end
          for (forvar238 = (1'h0); (forvar238 < (2'h3)); forvar238 = (forvar238 + (1'h1)))
            begin
              reg239 <= $unsigned(forvar106);
              reg240 = (((^((forvar195 ? wire229 : (8'hb4)) ?
                          (~reg180) : (reg211 ? reg133 : reg147))) ?
                      ((~$signed((8'ha5))) ?
                          (^reg107) : ($signed(reg161) ?
                              reg138 : $unsigned(reg220))) : forvar201[(3'h4):(1'h1)]) ?
                  reg218[(1'h0):(1'h0)] : ((($unsigned(forvar238) ^ ((8'hb1) + reg98)) ?
                      $unsigned({reg90}) : ($signed(forvar123) * reg213)) ^~ $signed(((reg94 ?
                          (8'h9f) : (8'ha5)) ?
                      {reg215} : reg207[(4'hb):(3'h6)]))));
              reg241 <= $unsigned({($unsigned(reg184) | reg93)});
              reg242 = $unsigned(reg162[(3'h7):(2'h3)]);
              reg243 <= reg127[(2'h2):(1'h0)];
            end
          for (forvar244 = (1'h0); (forvar244 < (2'h2)); forvar244 = (forvar244 + (1'h1)))
            begin
              reg245 = forvar244[(4'ha):(1'h0)];
              reg246 <= "QuQNEE";
              reg247 <= (reg199[(1'h1):(1'h1)] ? reg121 : reg216);
              reg248 <= (~(&{$signed((reg95 ? reg242 : forvar195)),
                  forvar186}));
            end
          reg249 <= $unsigned((({(reg143 & reg184), reg104[(1'h1):(1'h0)]} ?
                  (8'ha9) : $signed(forvar148[(2'h2):(1'h1)])) ?
              (((reg235 ? wire83 : reg245) ? reg146 : {reg219}) ?
                  (^(reg206 ?
                      reg134 : (7'h41))) : (((8'hb0) ^ reg89) << (&reg206))) : reg241));
        end
    end
  assign wire250 = (!(8'ha6));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1003
#( parameter param1132 = ({(((8'had) ? (^~(7'h43)) : ((7'h42) > (8'hbc))) <= {(~|(8'hb9))})} ? {(~|(((7'h40) | (8'h9f)) ? ((8'hb3) >>> (8'ha0)) : ((8'hbc) > (7'h40)))), ((^(8'hbf)) && (((8'ha5) ? (8'hb8) : (8'hac)) ? {(8'hab), (8'hb8)} : (&(8'ha9))))} : (|((-((8'hbe) ? (8'hab) : (8'hb5))) - (&{(8'hb1)}))))
, parameter param1133 = (~(((param1132 != {param1132, param1132}) ? param1132 : param1132) ? (&(param1132 ? param1132 : (param1132 <<< param1132))) : ((param1132 ? {param1132, param1132} : (param1132 ? param1132 : (7'h44))) << ((~(8'had)) & (param1132 ? param1132 : param1132))))) )
(y, clk, wire1008, wire1007, wire1006, wire1005, wire1004);
  output wire [(32'h59f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire1008;
  input wire signed [(4'h9):(1'h0)] wire1007;
  input wire [(5'h12):(1'h0)] wire1006;
  input wire [(4'hb):(1'h0)] wire1005;
  input wire signed [(2'h3):(1'h0)] wire1004;
  reg [(4'hf):(1'h0)] reg1131 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1130 = (1'h0);
  reg [(5'h14):(1'h0)] reg1129 = (1'h0);
  reg [(5'h15):(1'h0)] reg1128 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1127 = (1'h0);
  reg [(3'h4):(1'h0)] reg1126 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1125 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar1124 = (1'h0);
  reg [(2'h3):(1'h0)] reg1123 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire1122;
  wire [(5'h13):(1'h0)] wire1121;
  wire signed [(3'h5):(1'h0)] wire1120;
  reg [(2'h3):(1'h0)] reg1119 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1118 = (1'h0);
  reg [(4'ha):(1'h0)] reg1117 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1116 = (1'h0);
  reg [(3'h4):(1'h0)] reg1115 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1114 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1113 = (1'h0);
  reg [(2'h2):(1'h0)] reg1112 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1111 = (1'h0);
  reg [(5'h12):(1'h0)] reg1110 = (1'h0);
  reg [(5'h12):(1'h0)] reg1109 = (1'h0);
  reg [(5'h15):(1'h0)] reg1108 = (1'h0);
  reg [(4'ha):(1'h0)] reg1107 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1106 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1105 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1104 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1103 = (1'h0);
  wire [(2'h2):(1'h0)] wire1102;
  reg [(3'h5):(1'h0)] reg1101 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1100 = (1'h0);
  reg [(5'h12):(1'h0)] reg1099 = (1'h0);
  reg [(5'h14):(1'h0)] reg1098 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1097 = (1'h0);
  reg [(4'hd):(1'h0)] reg1096 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1095 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1094 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1093 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1092 = (1'h0);
  reg [(2'h2):(1'h0)] reg1091 = (1'h0);
  reg [(2'h3):(1'h0)] reg1084 = (1'h0);
  reg [(4'he):(1'h0)] reg1090 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1089 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1088 = (1'h0);
  reg [(5'h14):(1'h0)] reg1087 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1086 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1085 = (1'h0);
  reg [(4'he):(1'h0)] forvar1084 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1083 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1082 = (1'h0);
  reg [(4'ha):(1'h0)] reg1081 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1080 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1079 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1078 = (1'h0);
  wire signed [(2'h2):(1'h0)] wire1077;
  wire [(2'h3):(1'h0)] wire1076;
  reg [(4'h8):(1'h0)] reg1075 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1074 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1073 = (1'h0);
  reg [(5'h12):(1'h0)] reg1072 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1071 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1070 = (1'h0);
  reg [(3'h5):(1'h0)] reg1069 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1068 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1067 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1066 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1065 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1064 = (1'h0);
  reg [(3'h5):(1'h0)] reg1063 = (1'h0);
  reg [(3'h5):(1'h0)] reg1062 = (1'h0);
  reg [(4'h8):(1'h0)] reg1061 = (1'h0);
  reg [(2'h3):(1'h0)] reg1060 = (1'h0);
  reg [(4'h8):(1'h0)] reg1059 = (1'h0);
  reg [(5'h11):(1'h0)] reg1058 = (1'h0);
  wire signed [(5'h14):(1'h0)] wire1057;
  reg signed [(2'h3):(1'h0)] reg1049 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1043 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1042 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1056 = (1'h0);
  reg [(5'h13):(1'h0)] reg1055 = (1'h0);
  reg [(4'h8):(1'h0)] reg1054 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1053 = (1'h0);
  reg [(5'h13):(1'h0)] reg1052 = (1'h0);
  reg [(3'h6):(1'h0)] reg1051 = (1'h0);
  reg [(4'ha):(1'h0)] reg1050 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1049 = (1'h0);
  reg [(2'h2):(1'h0)] reg1048 = (1'h0);
  reg [(3'h5):(1'h0)] reg1047 = (1'h0);
  reg [(5'h15):(1'h0)] reg1046 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1045 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1044 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1043 = (1'h0);
  reg [(4'hf):(1'h0)] reg1042 = (1'h0);
  wire [(5'h12):(1'h0)] wire1041;
  wire signed [(3'h7):(1'h0)] wire1040;
  reg signed [(4'ha):(1'h0)] reg1031 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1030 = (1'h0);
  reg [(5'h14):(1'h0)] reg1039 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1038 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1037 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1036 = (1'h0);
  reg [(3'h4):(1'h0)] reg1035 = (1'h0);
  reg [(4'h9):(1'h0)] reg1034 = (1'h0);
  reg [(3'h7):(1'h0)] reg1033 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1032 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1031 = (1'h0);
  reg [(4'hb):(1'h0)] reg1030 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1029 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1028 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1027 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1026 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1025 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1024 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1023 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1022 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1021 = (1'h0);
  reg [(5'h10):(1'h0)] reg1020 = (1'h0);
  reg [(3'h7):(1'h0)] reg1019 = (1'h0);
  reg [(4'hb):(1'h0)] reg1018 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1014 = (1'h0);
  reg [(4'hb):(1'h0)] reg1012 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1017 = (1'h0);
  reg [(3'h4):(1'h0)] reg1016 = (1'h0);
  reg [(4'he):(1'h0)] reg1015 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1014 = (1'h0);
  reg [(3'h4):(1'h0)] reg1013 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1012 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1011 = (1'h0);
  wire [(4'hc):(1'h0)] wire1010;
  wire signed [(4'he):(1'h0)] wire1009;
  assign y = {reg1131,
                 reg1130,
                 reg1129,
                 reg1128,
                 forvar1127,
                 reg1126,
                 forvar1125,
                 forvar1124,
                 reg1123,
                 wire1122,
                 wire1121,
                 wire1120,
                 reg1119,
                 reg1118,
                 reg1117,
                 forvar1116,
                 reg1115,
                 reg1114,
                 reg1113,
                 reg1112,
                 forvar1111,
                 reg1110,
                 reg1109,
                 reg1108,
                 reg1107,
                 reg1106,
                 forvar1105,
                 reg1104,
                 forvar1103,
                 wire1102,
                 reg1101,
                 reg1100,
                 reg1099,
                 reg1098,
                 forvar1097,
                 reg1096,
                 reg1095,
                 reg1094,
                 forvar1093,
                 forvar1092,
                 reg1091,
                 reg1084,
                 reg1090,
                 reg1089,
                 reg1088,
                 reg1087,
                 reg1086,
                 reg1085,
                 forvar1084,
                 reg1083,
                 reg1082,
                 reg1081,
                 reg1080,
                 forvar1079,
                 reg1078,
                 wire1077,
                 wire1076,
                 reg1075,
                 reg1074,
                 forvar1073,
                 reg1072,
                 forvar1071,
                 reg1070,
                 reg1069,
                 forvar1068,
                 forvar1067,
                 reg1066,
                 reg1065,
                 reg1064,
                 reg1063,
                 reg1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 wire1057,
                 reg1049,
                 reg1043,
                 forvar1042,
                 reg1056,
                 reg1055,
                 reg1054,
                 forvar1053,
                 reg1052,
                 reg1051,
                 reg1050,
                 forvar1049,
                 reg1048,
                 reg1047,
                 reg1046,
                 reg1045,
                 reg1044,
                 forvar1043,
                 reg1042,
                 wire1041,
                 wire1040,
                 reg1031,
                 forvar1030,
                 reg1039,
                 reg1038,
                 forvar1037,
                 reg1036,
                 reg1035,
                 reg1034,
                 reg1033,
                 reg1032,
                 forvar1031,
                 reg1030,
                 reg1029,
                 reg1028,
                 reg1027,
                 reg1026,
                 reg1025,
                 reg1024,
                 forvar1023,
                 forvar1022,
                 reg1021,
                 reg1020,
                 reg1019,
                 reg1018,
                 reg1014,
                 reg1012,
                 reg1017,
                 reg1016,
                 reg1015,
                 forvar1014,
                 reg1013,
                 forvar1012,
                 reg1011,
                 wire1010,
                 wire1009,
                 (1'h0)};
  assign wire1009 = wire1007;
  assign wire1010 = ({wire1009[(4'h9):(4'h8)]} ?
                        (~&(wire1008[(1'h0):(1'h0)] ?
                            $signed((wire1007 || wire1009)) : (+wire1006))) : $signed(wire1004[(1'h0):(1'h0)]));
  always
    @(posedge clk) begin
      reg1011 <= wire1007;
      if ({(wire1007[(3'h4):(1'h1)] ?
              wire1006[(3'h4):(1'h1)] : ((|((8'ha7) ?
                  wire1008 : (8'ha1))) >> ($unsigned(wire1005) & {wire1009})))})
        begin
          for (forvar1012 = (1'h0); (forvar1012 < (2'h3)); forvar1012 = (forvar1012 + (1'h1)))
            begin
              reg1013 <= $signed((wire1006[(3'h7):(1'h1)] ?
                  forvar1012[(4'h9):(2'h3)] : (({reg1011, wire1008} ?
                          forvar1012[(3'h5):(2'h2)] : (wire1009 ?
                              wire1006 : wire1009)) ?
                      $unsigned((wire1004 ? (8'ha9) : wire1008)) : wire1008)));
            end
          for (forvar1014 = (1'h0); (forvar1014 < (3'h4)); forvar1014 = (forvar1014 + (1'h1)))
            begin
              reg1015 <= $unsigned($signed((wire1007[(3'h5):(1'h1)] ?
                  $signed(wire1009[(3'h5):(3'h5)]) : (wire1008 ?
                      reg1011[(2'h3):(2'h3)] : (&reg1013)))));
              reg1016 <= (reg1011 ^ (wire1010 >= $signed($unsigned($unsigned(wire1009)))));
            end
          reg1017 <= $unsigned($unsigned(wire1009));
        end
      else
        begin
          reg1012 = reg1017;
          if ($unsigned(((7'h43) == $signed($signed((reg1015 == reg1011))))))
            begin
              reg1013 = forvar1014;
              reg1014 = wire1010[(3'h7):(3'h6)];
              reg1015 = ($signed($unsigned(forvar1014)) ?
                  wire1006[(2'h3):(1'h0)] : wire1009);
              reg1016 = wire1007;
            end
          else
            begin
              reg1013 = $unsigned({$unsigned((~&$unsigned(forvar1012)))});
              reg1014 = {forvar1012};
              reg1015 <= {wire1008[(1'h0):(1'h0)],
                  ($unsigned(forvar1012) ?
                      $signed(({reg1017,
                          wire1010} ^~ $unsigned(forvar1012))) : (!$unsigned(wire1004[(1'h1):(1'h1)])))};
              reg1016 <= reg1015;
              reg1017 = wire1006[(5'h12):(3'h4)];
            end
          if (($unsigned((~(|$unsigned(wire1004)))) ?
              $signed((^wire1007[(3'h4):(2'h2)])) : reg1016[(3'h4):(2'h2)]))
            begin
              reg1018 <= reg1017[(1'h0):(1'h0)];
              reg1019 <= (&(-((~|$unsigned(wire1009)) ?
                  (|$signed(reg1011)) : wire1006[(4'hc):(4'hc)])));
              reg1020 <= forvar1012;
            end
          else
            begin
              reg1018 = (($unsigned((reg1016 ?
                          $unsigned((8'hb2)) : (wire1005 >>> reg1012))) ?
                      (8'h9f) : $signed(forvar1012[(5'h10):(3'h6)])) ?
                  reg1014 : (~(7'h44)));
              reg1019 <= reg1018;
            end
        end
      reg1021 <= wire1008;
    end
  always
    @(posedge clk) begin
      for (forvar1022 = (1'h0); (forvar1022 < (1'h0)); forvar1022 = (forvar1022 + (1'h1)))
        begin
          for (forvar1023 = (1'h0); (forvar1023 < (1'h1)); forvar1023 = (forvar1023 + (1'h1)))
            begin
              reg1024 <= (^$unsigned(({reg1020,
                      (reg1019 ? forvar1023 : wire1006)} ?
                  reg1018[(1'h0):(1'h0)] : forvar1014[(4'hb):(4'h9)])));
              reg1025 <= $unsigned($signed(((wire1004[(2'h3):(2'h3)] ?
                      ((7'h41) || wire1005) : $signed(reg1020)) ?
                  $unsigned((&reg1020)) : (+reg1011[(2'h2):(1'h1)]))));
              reg1026 = ((reg1011[(1'h1):(1'h0)] == $unsigned($unsigned(reg1025))) ?
                  forvar1023[(4'hd):(1'h0)] : $signed(({$signed((8'hae))} < wire1009[(3'h6):(3'h6)])));
              reg1027 = reg1014;
              reg1028 <= (8'had);
            end
          reg1029 <= (~wire1010[(4'ha):(4'ha)]);
        end
      if (wire1010[(4'hc):(3'h5)])
        begin
          reg1030 <= (reg1029[(1'h1):(1'h1)] ?
              {reg1014, $signed(reg1029)} : reg1028);
          for (forvar1031 = (1'h0); (forvar1031 < (1'h0)); forvar1031 = (forvar1031 + (1'h1)))
            begin
              reg1032 <= $unsigned((^(!({reg1024} > $signed(reg1020)))));
              reg1033 = (!("Vxx70r3EpwX" ?
                  ("lUiYq9" == $signed((^~reg1019))) : $unsigned(reg1025[(1'h0):(1'h0)])));
              reg1034 = ((^~(((~reg1025) * (forvar1023 ?
                      reg1018 : wire1005)) >= ((+wire1004) < $signed(forvar1031)))) ?
                  $unsigned((~|(&$unsigned((8'ha2))))) : ({reg1027[(4'h9):(1'h0)]} ?
                      (reg1032 ^ $unsigned(reg1029[(2'h3):(2'h3)])) : $unsigned(((wire1005 ?
                          reg1021 : forvar1031) >> $unsigned(forvar1031)))));
            end
          reg1035 <= {reg1026,
              ((!$unsigned(reg1033[(1'h1):(1'h1)])) ?
                  $unsigned($unsigned(((8'haa) ?
                      reg1015 : forvar1022))) : reg1013[(3'h4):(3'h4)])};
          reg1036 <= $unsigned((((7'h44) || forvar1023[(4'h9):(4'h8)]) - ($unsigned(((8'h9c) ?
                  wire1009 : reg1029)) ?
              $unsigned({wire1008}) : $signed($unsigned((8'ha8))))));
          for (forvar1037 = (1'h0); (forvar1037 < (2'h3)); forvar1037 = (forvar1037 + (1'h1)))
            begin
              reg1038 <= reg1030[(3'h4):(1'h0)];
              reg1039 <= $signed((reg1029 ?
                  forvar1031[(3'h4):(3'h4)] : ($signed((reg1033 ?
                          forvar1022 : (8'ha7))) ?
                      ((reg1032 ~^ reg1026) << {forvar1012,
                          reg1026}) : forvar1023[(4'hf):(4'ha)])));
            end
        end
      else
        begin
          for (forvar1030 = (1'h0); (forvar1030 < (1'h1)); forvar1030 = (forvar1030 + (1'h1)))
            begin
              reg1031 <= (reg1034 <= $signed(forvar1012[(4'h9):(1'h0)]));
              reg1032 <= (~|(8'hbb));
              reg1033 <= {$signed($signed($signed(reg1021)))};
            end
          reg1034 = (~|{forvar1023, "PkxOtq"});
        end
    end
  assign wire1040 = reg1015;
  assign wire1041 = ((forvar1022[(1'h0):(1'h0)] ~^ $unsigned(wire1010)) ?
                        {$unsigned($unsigned((~^reg1034)))} : (((~|{reg1011}) < ((8'ha2) <<< $signed(reg1012))) ?
                            {(reg1032[(4'h9):(1'h1)] ?
                                    wire1007[(1'h1):(1'h0)] : (forvar1037 | reg1029))} : {{$unsigned(reg1038),
                                    reg1031},
                                (forvar1031[(3'h6):(1'h1)] > forvar1014)}));
  always
    @(posedge clk) begin
      if ($unsigned((reg1011 ?
          $unsigned((reg1028 >>> ((8'hbe) | (8'ha2)))) : {($unsigned(reg1016) ^~ $unsigned(reg1039))})))
        begin
          reg1042 <= $signed((reg1030 ?
              ({$signed((8'hba)), ((8'hab) ? reg1033 : (8'ha5))} ?
                  (!(forvar1022 ? wire1006 : wire1040)) : {wire1005,
                      (+reg1029)}) : $signed((-"WP37HG2osAtkLMsyPgXk"))));
          for (forvar1043 = (1'h0); (forvar1043 < (2'h3)); forvar1043 = (forvar1043 + (1'h1)))
            begin
              reg1044 <= reg1021[(2'h3):(1'h0)];
              reg1045 <= $signed((&(forvar1030 ?
                  (forvar1030[(2'h2):(1'h0)] ^ reg1036) : ({reg1015} ?
                      (+forvar1022) : "0464qwT"))));
              reg1046 = (reg1015[(4'he):(4'hb)] != reg1012[(1'h1):(1'h0)]);
              reg1047 <= $unsigned(reg1033);
              reg1048 = ((+($signed((wire1006 * reg1015)) ?
                  $unsigned((reg1028 ~^ wire1040)) : ((wire1006 >> reg1034) ?
                      reg1045 : $signed(wire1006)))) >= $signed(reg1027));
            end
          for (forvar1049 = (1'h0); (forvar1049 < (3'h4)); forvar1049 = (forvar1049 + (1'h1)))
            begin
              reg1050 <= $unsigned("iwnKYIDIrRSnv");
              reg1051 <= (forvar1037[(1'h1):(1'h0)] ?
                  (reg1029 ^ {reg1039[(5'h10):(4'hd)]}) : (^~reg1030));
              reg1052 <= (!$signed($unsigned($unsigned((wire1040 > reg1050)))));
            end
          for (forvar1053 = (1'h0); (forvar1053 < (2'h2)); forvar1053 = (forvar1053 + (1'h1)))
            begin
              reg1054 = $unsigned(forvar1043[(3'h7):(3'h6)]);
              reg1055 = reg1046[(3'h7):(1'h0)];
              reg1056 = (~((forvar1012 ?
                  (~^(-forvar1043)) : {{reg1017, reg1015},
                      reg1036[(1'h1):(1'h0)]}) > reg1015));
            end
        end
      else
        begin
          for (forvar1042 = (1'h0); (forvar1042 < (1'h0)); forvar1042 = (forvar1042 + (1'h1)))
            begin
              reg1043 = reg1055;
              reg1044 = (-reg1052[(4'ha):(4'ha)]);
              reg1045 = "0BHHzZNqY0JilI";
              reg1046 = $signed(($signed((-$unsigned(reg1024))) > $signed((!(wire1007 ?
                  (7'h44) : wire1040)))));
            end
          if ($signed((8'ha4)))
            begin
              reg1047 <= $signed(wire1008[(1'h1):(1'h0)]);
              reg1048 <= ((reg1036 ?
                      $signed($unsigned(reg1024)) : ((reg1052[(4'hc):(3'h5)] ?
                          reg1019[(3'h4):(2'h3)] : "y0sU") + $signed(reg1045[(3'h5):(1'h0)]))) ?
                  $unsigned(((^$signed((8'ha7))) ?
                      $unsigned((reg1029 ^~ wire1006)) : {$unsigned(reg1012)})) : ($unsigned((((8'ha8) - reg1019) <= ((8'ha6) ?
                      forvar1031 : reg1036))) & reg1032));
              reg1049 = reg1029;
              reg1050 <= $signed(((($unsigned((8'h9c)) ?
                  reg1052 : (-forvar1014)) >= ($signed(reg1031) ?
                  $signed(wire1010) : $unsigned(reg1034))) || (+$unsigned({reg1030,
                  wire1004}))));
            end
          else
            begin
              reg1047 = {$signed($signed((forvar1031 != "v"))),
                  ($unsigned(((reg1018 ?
                      forvar1023 : reg1050) ^~ $unsigned(reg1055))) >>> ((wire1041[(4'h8):(3'h4)] ?
                          $unsigned(reg1017) : $signed(reg1039)) ?
                      $signed($signed(reg1031)) : wire1040[(3'h4):(2'h3)]))};
              reg1048 = reg1046[(3'h7):(3'h7)];
            end
        end
    end
  assign wire1057 = ($signed(forvar1023) ?
                        reg1015 : ((|reg1033) ?
                            $signed(($signed((8'ha3)) || (reg1027 ~^ reg1036))) : "HG"));
  always
    @(posedge clk) begin
      if ($signed($signed($unsigned(reg1033))))
        begin
          reg1058 <= ((&$signed({reg1044[(3'h4):(3'h4)],
              (8'hbc)})) ~^ {(~$unsigned((|wire1004)))});
          reg1059 = reg1016;
          if (reg1059[(2'h3):(1'h0)])
            begin
              reg1060 = $signed((~|($signed($unsigned((8'h9e))) < ((wire1006 ?
                      reg1029 : forvar1030) ?
                  reg1038 : {reg1030}))));
              reg1061 = {(({(8'ha6)} << reg1026[(5'h12):(4'hc)]) | ($signed((~forvar1049)) ?
                      (~$unsigned((8'hbb))) : (^~reg1049[(2'h2):(1'h0)]))),
                  (reg1024[(3'h4):(2'h2)] ?
                      reg1032 : ($signed($unsigned(wire1008)) == $signed($signed(reg1052))))};
              reg1062 = reg1027[(3'h7):(3'h5)];
              reg1063 = {forvar1022};
              reg1064 = $unsigned($unsigned(reg1032[(2'h2):(1'h1)]));
            end
          else
            begin
              reg1060 <= (reg1021 >= ((~|forvar1030) && wire1041[(2'h2):(2'h2)]));
              reg1061 <= reg1020;
              reg1062 <= ((($unsigned(wire1057[(3'h4):(1'h0)]) || reg1028[(3'h5):(3'h4)]) ?
                  wire1007[(3'h5):(3'h5)] : $signed($signed((reg1043 <<< reg1045)))) >= ($signed($unsigned($unsigned(forvar1037))) ?
                  $unsigned(reg1034) : (reg1039[(4'hf):(1'h1)] ?
                      reg1035 : $signed($unsigned(reg1064)))));
              reg1063 <= (~($signed(wire1040) << $unsigned("VMveBNXvBYV")));
              reg1064 = $unsigned(reg1030);
            end
          reg1065 = $signed((({reg1015[(3'h7):(2'h3)], (+forvar1014)} ?
              ((forvar1031 ?
                  wire1040 : reg1060) - reg1062) : reg1046[(3'h5):(1'h0)]) << (reg1055[(4'hd):(3'h7)] <<< (reg1062[(3'h4):(2'h2)] ?
              (reg1031 & reg1048) : reg1059[(1'h1):(1'h0)]))));
          reg1066 <= ($unsigned($signed(reg1060[(2'h3):(2'h3)])) ?
              reg1029 : reg1047[(1'h1):(1'h1)]);
        end
      else
        begin
          reg1058 <= ((~^(($signed(reg1024) <<< "5HIvpBXvlXsAam86F4") >= (&{reg1020}))) ?
              $unsigned(reg1063) : (&reg1047[(1'h1):(1'h1)]));
          if ($unsigned(($signed(reg1055[(4'hc):(2'h3)]) ?
              ($unsigned(reg1029) ? reg1011 : reg1038) : (forvar1012 ?
                  ("5GQiD5" ^ (reg1021 ^~ reg1031)) : ($unsigned(reg1034) != (reg1065 >>> (7'h43)))))))
            begin
              reg1059 <= (&(wire1005 ?
                  {"Hn1t"} : (|$unsigned("urDunxtzd53wb"))));
              reg1060 <= $unsigned($unsigned((|$signed((!forvar1022)))));
              reg1061 <= reg1020[(4'hb):(3'h4)];
              reg1062 <= reg1052;
            end
          else
            begin
              reg1059 = ((reg1017[(1'h1):(1'h0)] ?
                  ($signed((wire1006 ?
                      reg1031 : reg1062)) <<< (~"UbYoMKmPKsnGHhmkUd")) : (|reg1051)) ^~ ($signed(reg1012[(1'h1):(1'h1)]) ?
                  reg1056 : reg1031));
              reg1060 <= $signed(reg1024[(1'h1):(1'h0)]);
              reg1061 <= reg1029;
              reg1062 <= reg1056[(4'hf):(3'h4)];
            end
        end
      for (forvar1067 = (1'h0); (forvar1067 < (1'h1)); forvar1067 = (forvar1067 + (1'h1)))
        begin
          for (forvar1068 = (1'h0); (forvar1068 < (1'h1)); forvar1068 = (forvar1068 + (1'h1)))
            begin
              reg1069 = (8'ha0);
              reg1070 <= $signed((reg1020[(4'hb):(4'h8)] ?
                  (reg1034[(4'h8):(4'h8)] - $signed((forvar1053 + reg1049))) : ($unsigned((~&reg1048)) <= $signed($unsigned(reg1033)))));
            end
        end
      for (forvar1071 = (1'h0); (forvar1071 < (2'h3)); forvar1071 = (forvar1071 + (1'h1)))
        begin
          reg1072 = wire1008[(1'h0):(1'h0)];
          for (forvar1073 = (1'h0); (forvar1073 < (1'h0)); forvar1073 = (forvar1073 + (1'h1)))
            begin
              reg1074 = forvar1014[(3'h6):(1'h1)];
            end
          reg1075 <= (forvar1049[(3'h5):(1'h0)] ?
              (~^($unsigned((reg1061 ? reg1056 : reg1043)) ?
                  (|$unsigned((8'hb5))) : forvar1067)) : wire1040[(3'h4):(1'h0)]);
        end
    end
  assign wire1076 = reg1049[(1'h0):(1'h0)];
  assign wire1077 = reg1014[(3'h4):(2'h2)];
  always
    @(posedge clk) begin
      reg1078 = $signed($signed($signed($signed((8'h9f)))));
      if (reg1043)
        begin
          for (forvar1079 = (1'h0); (forvar1079 < (1'h1)); forvar1079 = (forvar1079 + (1'h1)))
            begin
              reg1080 <= ($unsigned(($unsigned({reg1065}) ?
                  wire1005 : {$unsigned(reg1069),
                      $signed(reg1050)})) >> $signed(forvar1071));
              reg1081 <= {(-$unsigned(wire1009[(4'he):(4'he)]))};
              reg1082 <= reg1016;
            end
          reg1083 = {$signed(reg1027[(4'hc):(2'h2)]),
              ((!$unsigned(wire1040[(2'h2):(1'h1)])) | reg1050)};
          for (forvar1084 = (1'h0); (forvar1084 < (2'h2)); forvar1084 = (forvar1084 + (1'h1)))
            begin
              reg1085 = (reg1011 - forvar1049[(3'h4):(1'h0)]);
              reg1086 = $signed(forvar1037);
              reg1087 <= reg1012[(3'h6):(3'h5)];
              reg1088 = $unsigned(($unsigned($signed($signed(reg1018))) ?
                  ({$unsigned(reg1020), (-wire1004)} ?
                      ((~^forvar1030) ?
                          reg1012 : (reg1085 ?
                              reg1087 : (8'had))) : $unsigned(reg1025)) : forvar1012[(4'ha):(4'ha)]));
              reg1089 <= forvar1068;
            end
          reg1090 <= ($signed(({$signed(reg1031)} ?
              (~|forvar1042) : $unsigned((8'ha2)))) - $unsigned("fDBV"));
        end
      else
        begin
          for (forvar1079 = (1'h0); (forvar1079 < (2'h3)); forvar1079 = (forvar1079 + (1'h1)))
            begin
              reg1080 <= reg1015;
              reg1081 <= forvar1037;
              reg1082 <= (~|(+(($unsigned(forvar1071) ?
                  (reg1088 ?
                      reg1042 : reg1028) : $signed(forvar1053)) ^~ ((reg1015 >= reg1013) ?
                  $signed(reg1064) : ((8'hae) ? reg1089 : (8'hac))))));
              reg1083 = $signed((&reg1066));
              reg1084 = (~|(^~{(~^(^~reg1074))}));
            end
        end
      reg1091 = reg1042;
      for (forvar1092 = (1'h0); (forvar1092 < (3'h4)); forvar1092 = (forvar1092 + (1'h1)))
        begin
          for (forvar1093 = (1'h0); (forvar1093 < (1'h0)); forvar1093 = (forvar1093 + (1'h1)))
            begin
              reg1094 <= forvar1022;
              reg1095 = $signed($unsigned(((+{(8'h9f)}) ?
                  $unsigned((reg1035 >>> reg1035)) : reg1014[(1'h1):(1'h0)])));
              reg1096 <= forvar1084;
            end
          for (forvar1097 = (1'h0); (forvar1097 < (1'h0)); forvar1097 = (forvar1097 + (1'h1)))
            begin
              reg1098 = (~(~|reg1038[(4'hc):(4'h8)]));
              reg1099 = $signed(reg1036);
              reg1100 <= forvar1071;
            end
        end
      reg1101 <= $unsigned(($unsigned(forvar1043) ? (+reg1051) : forvar1093));
    end
  assign wire1102 = reg1033;
  always
    @(posedge clk) begin
      for (forvar1103 = (1'h0); (forvar1103 < (3'h4)); forvar1103 = (forvar1103 + (1'h1)))
        begin
          reg1104 = "qdC7BDxKY7UEcCKmO9";
          for (forvar1105 = (1'h0); (forvar1105 < (1'h0)); forvar1105 = (forvar1105 + (1'h1)))
            begin
              reg1106 <= (|"QxM");
              reg1107 = reg1078;
              reg1108 <= $signed(forvar1023[(3'h4):(1'h1)]);
              reg1109 <= ((~&$unsigned(({reg1074} != $unsigned(reg1086)))) & reg1060[(1'h1):(1'h0)]);
              reg1110 <= {(forvar1068 > (+$signed($unsigned(reg1020))))};
            end
          for (forvar1111 = (1'h0); (forvar1111 < (2'h3)); forvar1111 = (forvar1111 + (1'h1)))
            begin
              reg1112 <= "anf1UiLIZlKSTVgdNcKd";
              reg1113 <= reg1069[(1'h1):(1'h1)];
              reg1114 = (forvar1031 + ((reg1014[(3'h5):(1'h1)] - $unsigned((reg1094 ^~ forvar1103))) ?
                  (|({forvar1042} ?
                      $signed(reg1069) : (reg1066 ?
                          reg1110 : reg1086))) : ($signed($unsigned(reg1098)) + (&$unsigned((8'hb3))))));
            end
          reg1115 = (7'h41);
          for (forvar1116 = (1'h0); (forvar1116 < (1'h0)); forvar1116 = (forvar1116 + (1'h1)))
            begin
              reg1117 <= (wire1008 ?
                  $signed($signed(((&reg1106) ?
                      $unsigned((8'hbd)) : reg1013[(2'h2):(1'h0)]))) : reg1016[(3'h4):(2'h3)]);
              reg1118 <= (8'hb9);
              reg1119 <= (reg1047[(1'h0):(1'h0)] ?
                  $unsigned((8'hb5)) : ("RDimJY1XNl" ?
                      ($unsigned((reg1060 >>> forvar1031)) ?
                          (!$unsigned(forvar1105)) : {reg1029[(1'h1):(1'h0)]}) : forvar1067[(4'he):(4'ha)]));
            end
        end
    end
  assign wire1120 = ("" ?
                        (~^(reg1081[(3'h4):(2'h3)] + (^$unsigned(forvar1053)))) : $signed(reg1072));
  assign wire1121 = $signed((&$signed(((reg1029 <= reg1049) ?
                        wire1009[(3'h4):(2'h2)] : ((8'hb2) >= reg1080)))));
  assign wire1122 = (^(forvar1111 & (reg1108 ?
                        $unsigned(forvar1116) : (reg1059 > (reg1059 ?
                            reg1030 : reg1087)))));
  always
    @(posedge clk) begin
      reg1123 <= {$signed((^$signed((reg1035 <= wire1010)))),
          ($signed(({reg1014, forvar1049} ?
                  $unsigned(reg1089) : (reg1063 | reg1087))) ?
              ($signed((reg1088 ?
                  reg1113 : reg1089)) == {reg1088[(2'h3):(1'h1)]}) : $unsigned("VZoL8J0Vq"))};
      for (forvar1124 = (1'h0); (forvar1124 < (3'h4)); forvar1124 = (forvar1124 + (1'h1)))
        begin
          for (forvar1125 = (1'h0); (forvar1125 < (2'h2)); forvar1125 = (forvar1125 + (1'h1)))
            begin
              reg1126 <= $unsigned($unsigned($signed((|((8'h9d) < reg1011)))));
            end
          for (forvar1127 = (1'h0); (forvar1127 < (1'h1)); forvar1127 = (forvar1127 + (1'h1)))
            begin
              reg1128 <= reg1062[(3'h5):(3'h4)];
              reg1129 = ((reg1086[(4'hc):(2'h2)] >>> $unsigned($unsigned($signed(reg1118)))) || {($unsigned($unsigned(reg1115)) ?
                      (reg1062[(1'h1):(1'h1)] | (wire1009 ?
                          reg1082 : (8'hac))) : reg1052[(3'h6):(1'h0)]),
                  ({reg1064, (&reg1078)} >> $signed(reg1024))});
              reg1130 = ((~^$unsigned(reg1029)) ?
                  ((~|("y" ~^ (reg1118 && reg1110))) >>> {$unsigned($unsigned((8'ha2))),
                      (8'ha8)}) : ($signed(reg1106[(3'h4):(2'h2)]) != reg1014));
            end
          reg1131 = (!forvar1093[(4'hc):(4'hc)]);
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module818
#( parameter param997 = ({(!{(~(8'ha6)), {(7'h43), (7'h41)}})} && (((^~(~|(8'haf))) - ({(8'ha2)} << {(8'haa), (8'hac)})) ? ((!(!(8'ha3))) ? (((8'ha9) ? (8'ha4) : (8'ha0)) ? (&(8'had)) : ((8'h9c) ? (8'hb4) : (7'h44))) : (!((7'h43) < (8'hb4)))) : {(((8'haa) >> (8'hbd)) ? {(7'h41)} : (8'hbb))}))
, parameter param998 = (((({param997} ^ (^~param997)) ? param997 : param997) - param997) ? param997 : (~&(7'h44))) )
(y, clk, wire822, wire821, wire820, wire819);
  output wire [(32'h8cf):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire822;
  input wire [(4'ha):(1'h0)] wire821;
  input wire [(5'h11):(1'h0)] wire820;
  input wire signed [(4'ha):(1'h0)] wire819;
  reg signed [(4'he):(1'h0)] reg996 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg995 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg994 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar993 = (1'h0);
  reg [(4'h8):(1'h0)] reg992 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar991 = (1'h0);
  reg [(4'h9):(1'h0)] forvar990 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg989 = (1'h0);
  reg [(4'hf):(1'h0)] reg988 = (1'h0);
  reg [(5'h13):(1'h0)] reg987 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar986 = (1'h0);
  reg signed [(4'he):(1'h0)] reg985 = (1'h0);
  reg [(4'hf):(1'h0)] reg984 = (1'h0);
  reg [(4'he):(1'h0)] reg983 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg982 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg981 = (1'h0);
  reg [(5'h14):(1'h0)] reg980 = (1'h0);
  reg [(5'h13):(1'h0)] forvar979 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar978 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg977 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire976;
  reg [(5'h12):(1'h0)] reg975 = (1'h0);
  reg [(4'hc):(1'h0)] reg974 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar973 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg972 = (1'h0);
  reg [(4'hb):(1'h0)] reg971 = (1'h0);
  reg [(5'h10):(1'h0)] reg970 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg969 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg968 = (1'h0);
  reg [(3'h7):(1'h0)] forvar967 = (1'h0);
  reg [(4'hf):(1'h0)] reg966 = (1'h0);
  reg [(4'ha):(1'h0)] reg965 = (1'h0);
  reg [(3'h6):(1'h0)] forvar964 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg963 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar962 = (1'h0);
  reg [(5'h15):(1'h0)] reg961 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg960 = (1'h0);
  reg [(3'h6):(1'h0)] reg959 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg958 = (1'h0);
  reg [(4'he):(1'h0)] forvar957 = (1'h0);
  reg [(5'h12):(1'h0)] reg956 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg955 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg954 = (1'h0);
  reg signed [(4'he):(1'h0)] reg953 = (1'h0);
  reg [(3'h6):(1'h0)] forvar952 = (1'h0);
  reg [(4'h9):(1'h0)] forvar951 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg950 = (1'h0);
  reg [(2'h3):(1'h0)] reg949 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar948 = (1'h0);
  reg [(2'h2):(1'h0)] reg947 = (1'h0);
  reg [(3'h5):(1'h0)] reg946 = (1'h0);
  reg signed [(4'he):(1'h0)] reg945 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg944 = (1'h0);
  reg [(4'hb):(1'h0)] forvar943 = (1'h0);
  reg [(5'h12):(1'h0)] reg942 = (1'h0);
  reg [(4'hd):(1'h0)] reg941 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg940 = (1'h0);
  reg [(4'he):(1'h0)] forvar939 = (1'h0);
  reg [(3'h4):(1'h0)] reg938 = (1'h0);
  reg [(5'h11):(1'h0)] reg937 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar936 = (1'h0);
  reg [(3'h4):(1'h0)] reg935 = (1'h0);
  reg [(3'h6):(1'h0)] reg934 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg933 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg932 = (1'h0);
  reg [(2'h2):(1'h0)] reg931 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar930 = (1'h0);
  reg [(3'h6):(1'h0)] forvar929 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg928 = (1'h0);
  reg [(5'h15):(1'h0)] reg927 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg926 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg925 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg924 = (1'h0);
  reg [(2'h2):(1'h0)] reg923 = (1'h0);
  reg [(4'hb):(1'h0)] forvar922 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg922 = (1'h0);
  reg [(3'h6):(1'h0)] reg921 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg920 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg919 = (1'h0);
  reg signed [(4'he):(1'h0)] reg918 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg917 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg916 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar915 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg914 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg913 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg912 = (1'h0);
  reg [(5'h10):(1'h0)] reg911 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg910 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar909 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg908 = (1'h0);
  reg [(3'h5):(1'h0)] reg907 = (1'h0);
  reg [(4'ha):(1'h0)] reg906 = (1'h0);
  reg signed [(4'he):(1'h0)] reg905 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg904 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar903 = (1'h0);
  reg [(4'hf):(1'h0)] reg902 = (1'h0);
  reg [(5'h15):(1'h0)] reg901 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg899 = (1'h0);
  reg [(3'h5):(1'h0)] reg898 = (1'h0);
  reg [(5'h12):(1'h0)] forvar897 = (1'h0);
  wire [(5'h11):(1'h0)] wire896;
  wire signed [(4'h9):(1'h0)] wire895;
  wire [(4'ha):(1'h0)] wire894;
  wire [(4'he):(1'h0)] wire893;
  wire [(4'ha):(1'h0)] wire892;
  wire signed [(4'hb):(1'h0)] wire891;
  wire signed [(4'hc):(1'h0)] wire890;
  wire [(4'hc):(1'h0)] wire889;
  reg [(4'hc):(1'h0)] reg888 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg887 = (1'h0);
  reg [(4'he):(1'h0)] reg886 = (1'h0);
  reg [(5'h15):(1'h0)] reg885 = (1'h0);
  reg [(5'h10):(1'h0)] reg884 = (1'h0);
  reg [(4'ha):(1'h0)] reg883 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg882 = (1'h0);
  reg [(5'h11):(1'h0)] forvar881 = (1'h0);
  wire [(4'hd):(1'h0)] wire880;
  reg [(3'h6):(1'h0)] reg879 = (1'h0);
  reg [(2'h3):(1'h0)] reg878 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg877 = (1'h0);
  reg [(5'h10):(1'h0)] reg876 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg875 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg874 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg873 = (1'h0);
  reg [(2'h3):(1'h0)] forvar872 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg871 = (1'h0);
  reg [(4'hd):(1'h0)] reg870 = (1'h0);
  reg [(4'hd):(1'h0)] forvar869 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg868 = (1'h0);
  reg [(5'h14):(1'h0)] forvar867 = (1'h0);
  reg [(4'ha):(1'h0)] reg855 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg866 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg865 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg864 = (1'h0);
  reg [(4'he):(1'h0)] reg863 = (1'h0);
  reg [(5'h10):(1'h0)] reg862 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg861 = (1'h0);
  reg [(5'h12):(1'h0)] reg860 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg859 = (1'h0);
  reg signed [(4'he):(1'h0)] reg858 = (1'h0);
  reg [(4'ha):(1'h0)] reg857 = (1'h0);
  reg [(4'h8):(1'h0)] reg856 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar855 = (1'h0);
  reg [(5'h14):(1'h0)] reg854 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg853 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg852 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg850 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg849 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg848 = (1'h0);
  reg signed [(4'he):(1'h0)] reg847 = (1'h0);
  reg [(4'hd):(1'h0)] reg846 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg845 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg844 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar843 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar842 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg838 = (1'h0);
  reg [(4'hf):(1'h0)] forvar835 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg834 = (1'h0);
  reg [(4'hc):(1'h0)] forvar832 = (1'h0);
  reg [(2'h3):(1'h0)] reg831 = (1'h0);
  reg [(5'h14):(1'h0)] forvar829 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg827 = (1'h0);
  reg [(4'hb):(1'h0)] forvar826 = (1'h0);
  reg [(2'h3):(1'h0)] reg841 = (1'h0);
  reg [(4'hd):(1'h0)] reg840 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg839 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar838 = (1'h0);
  reg [(5'h13):(1'h0)] reg837 = (1'h0);
  reg [(5'h13):(1'h0)] reg836 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg835 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar834 = (1'h0);
  reg [(5'h13):(1'h0)] reg833 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg832 = (1'h0);
  reg [(4'h9):(1'h0)] forvar831 = (1'h0);
  reg [(5'h13):(1'h0)] reg830 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg829 = (1'h0);
  reg [(5'h10):(1'h0)] reg828 = (1'h0);
  reg [(4'h8):(1'h0)] forvar827 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg826 = (1'h0);
  wire signed [(5'h11):(1'h0)] wire825;
  wire signed [(4'he):(1'h0)] wire824;
  wire [(4'h8):(1'h0)] wire823;
  assign y = {reg996,
                 reg995,
                 reg994,
                 forvar993,
                 reg992,
                 forvar991,
                 forvar990,
                 reg989,
                 reg988,
                 reg987,
                 forvar986,
                 reg985,
                 reg984,
                 reg983,
                 reg982,
                 reg981,
                 reg980,
                 forvar979,
                 forvar978,
                 reg977,
                 wire976,
                 reg975,
                 reg974,
                 forvar973,
                 reg972,
                 reg971,
                 reg970,
                 reg969,
                 reg968,
                 forvar967,
                 reg966,
                 reg965,
                 forvar964,
                 reg963,
                 forvar962,
                 reg961,
                 reg960,
                 reg959,
                 reg958,
                 forvar957,
                 reg956,
                 reg955,
                 reg954,
                 reg953,
                 forvar952,
                 forvar951,
                 reg950,
                 reg949,
                 forvar948,
                 reg947,
                 reg946,
                 reg945,
                 reg944,
                 forvar943,
                 reg942,
                 reg941,
                 reg940,
                 forvar939,
                 reg938,
                 reg937,
                 forvar936,
                 reg935,
                 reg934,
                 reg933,
                 reg932,
                 reg931,
                 forvar930,
                 forvar929,
                 reg928,
                 reg927,
                 reg926,
                 reg925,
                 reg924,
                 reg923,
                 forvar922,
                 reg922,
                 reg921,
                 reg920,
                 reg919,
                 reg918,
                 reg917,
                 reg916,
                 forvar915,
                 reg914,
                 reg913,
                 reg912,
                 reg911,
                 reg910,
                 forvar909,
                 reg908,
                 reg907,
                 reg906,
                 reg905,
                 reg904,
                 forvar903,
                 reg902,
                 reg901,
                 reg900,
                 reg899,
                 reg898,
                 forvar897,
                 wire896,
                 wire895,
                 wire894,
                 wire893,
                 wire892,
                 wire891,
                 wire890,
                 wire889,
                 reg888,
                 reg887,
                 reg886,
                 reg885,
                 reg884,
                 reg883,
                 reg882,
                 forvar881,
                 wire880,
                 reg879,
                 reg878,
                 reg877,
                 reg876,
                 reg875,
                 reg874,
                 reg873,
                 forvar872,
                 reg871,
                 reg870,
                 forvar869,
                 reg868,
                 forvar867,
                 reg855,
                 reg866,
                 reg865,
                 reg864,
                 reg863,
                 reg862,
                 reg861,
                 reg860,
                 reg859,
                 reg858,
                 reg857,
                 reg856,
                 forvar855,
                 reg854,
                 reg853,
                 reg852,
                 reg851,
                 reg850,
                 reg849,
                 reg848,
                 reg847,
                 reg846,
                 reg845,
                 reg844,
                 forvar843,
                 forvar842,
                 reg838,
                 forvar835,
                 reg834,
                 forvar832,
                 reg831,
                 forvar829,
                 reg827,
                 forvar826,
                 reg841,
                 reg840,
                 reg839,
                 forvar838,
                 reg837,
                 reg836,
                 reg835,
                 forvar834,
                 reg833,
                 reg832,
                 forvar831,
                 reg830,
                 reg829,
                 reg828,
                 forvar827,
                 reg826,
                 wire825,
                 wire824,
                 wire823,
                 (1'h0)};
  assign wire823 = {(~wire820),
                       ((((wire820 ?
                               wire821 : (8'ha6)) ^~ (wire820 - wire822)) <= wire821[(3'h5):(1'h1)]) ?
                           wire821[(2'h2):(2'h2)] : $unsigned(wire821[(3'h4):(1'h0)]))};
  assign wire824 = wire819[(3'h4):(3'h4)];
  assign wire825 = (($signed($signed($signed(wire820))) ?
                       "BXsDVxlaZgmA6" : (~wire821)) >>> (+((8'hb1) ?
                       (~{wire822, wire820}) : (|((7'h41) ?
                           wire821 : wire823)))));
  always
    @(posedge clk) begin
      if ((wire824[(4'h8):(1'h1)] >= (wire821 | $signed($unsigned($signed(wire824))))))
        begin
          reg826 <= wire820;
          for (forvar827 = (1'h0); (forvar827 < (2'h3)); forvar827 = (forvar827 + (1'h1)))
            begin
              reg828 <= (~^{$unsigned(((wire821 <<< forvar827) || (wire822 & reg826)))});
              reg829 = (^($unsigned((~^(&wire824))) ?
                  (wire823[(4'h8):(3'h7)] - (-wire819)) : wire821));
              reg830 = "dhMcrQBO6f270bIgbo";
            end
          for (forvar831 = (1'h0); (forvar831 < (1'h1)); forvar831 = (forvar831 + (1'h1)))
            begin
              reg832 <= (^~(^({$unsigned(reg826)} >> "LPCcOdmU")));
              reg833 = (8'hba);
            end
          for (forvar834 = (1'h0); (forvar834 < (1'h0)); forvar834 = (forvar834 + (1'h1)))
            begin
              reg835 = $signed({"ELffTemPIBHq",
                  {reg829[(3'h4):(2'h2)], forvar834}});
              reg836 = (({$unsigned(reg830), (8'hb7)} ?
                  "d3l01iUHRnYgM" : reg835) == (reg826[(3'h4):(1'h1)] ?
                  wire823 : $unsigned(reg833[(4'h9):(3'h6)])));
              reg837 <= (8'haa);
            end
          for (forvar838 = (1'h0); (forvar838 < (2'h3)); forvar838 = (forvar838 + (1'h1)))
            begin
              reg839 <= (((reg830 ?
                  (+reg830) : ($signed(wire822) != {(8'ha3)})) >>> reg836[(3'h6):(3'h4)]) < $unsigned($unsigned((reg826[(4'h8):(3'h7)] > $signed((8'had))))));
              reg840 <= "AIpUWA6m4rIn";
              reg841 <= ({wire819, reg835} != $unsigned($signed({reg829})));
            end
        end
      else
        begin
          for (forvar826 = (1'h0); (forvar826 < (2'h2)); forvar826 = (forvar826 + (1'h1)))
            begin
              reg827 = $unsigned($unsigned($unsigned(reg840)));
              reg828 <= reg836[(3'h5):(1'h0)];
            end
          for (forvar829 = (1'h0); (forvar829 < (2'h2)); forvar829 = (forvar829 + (1'h1)))
            begin
              reg830 = wire819;
              reg831 = $unsigned($signed(reg835));
            end
          for (forvar832 = (1'h0); (forvar832 < (2'h3)); forvar832 = (forvar832 + (1'h1)))
            begin
              reg833 <= (((-(!$signed(reg828))) ?
                  ($unsigned((|wire820)) ?
                      wire821 : ($signed((8'h9e)) ?
                          (forvar829 < reg841) : reg833[(3'h7):(1'h1)])) : $unsigned($signed((forvar834 ?
                      forvar826 : reg841)))) && $unsigned(((-reg833) ~^ $signed((reg837 ?
                  forvar832 : forvar831)))));
              reg834 <= "PcaLCXsFr7sN";
            end
          for (forvar835 = (1'h0); (forvar835 < (1'h1)); forvar835 = (forvar835 + (1'h1)))
            begin
              reg836 <= (forvar827 ?
                  ((^((^~wire825) >> ((8'hb6) ?
                      reg831 : reg835))) | forvar831) : $unsigned({(-forvar826[(3'h5):(1'h0)])}));
              reg837 <= $signed(forvar835);
              reg838 <= reg835[(1'h1):(1'h1)];
            end
        end
      for (forvar842 = (1'h0); (forvar842 < (3'h4)); forvar842 = (forvar842 + (1'h1)))
        begin
          for (forvar843 = (1'h0); (forvar843 < (2'h2)); forvar843 = (forvar843 + (1'h1)))
            begin
              reg844 <= $signed($signed($unsigned((~&(~^forvar834)))));
            end
          if ((~(^~(wire822 ?
              $unsigned((forvar832 <= (8'hac))) : {{(8'ha2)},
                  (forvar829 ? forvar835 : wire820)}))))
            begin
              reg845 <= $unsigned(forvar826[(3'h7):(3'h5)]);
              reg846 = forvar829[(5'h10):(3'h7)];
              reg847 <= ((~(7'h40)) - ("DDXcmhS4" ~^ (^~reg841)));
              reg848 = "hVYFFB2whW";
              reg849 <= ($signed((((+forvar835) ?
                          wire825[(3'h7):(2'h2)] : $signed(reg830)) ?
                      ($signed(forvar829) ?
                          $signed((8'hb4)) : (reg847 ?
                              reg844 : wire825)) : ({reg834, reg839} ?
                          "G1xuwMalKVKm" : {forvar827}))) ?
                  (^(((^~(8'hbb)) ?
                          (reg848 ?
                              wire820 : forvar835) : reg832[(3'h5):(2'h3)]) ?
                      (((8'ha5) ^ reg845) != (reg845 ?
                          reg835 : (8'hae))) : (8'ha7))) : (^({{reg833}} ?
                      wire825[(4'he):(1'h0)] : (reg833 ?
                          (wire825 >= (8'hb8)) : $signed((8'haf))))));
            end
          else
            begin
              reg845 = ((wire823 + (~|(~(^reg841)))) ^~ $signed($signed(((reg826 ?
                  reg847 : wire823) <= reg830[(5'h10):(1'h1)]))));
              reg846 <= forvar829;
              reg847 = (((~(reg836[(5'h10):(4'ha)] & wire821)) ?
                      ({{forvar829, (7'h42)}} > reg849) : (reg846 ?
                          reg848 : ("B8Zxpyzqa54HmEVuu9" >>> {reg849}))) ?
                  $signed("rOI") : ((reg835 ?
                      ((&forvar834) || ((8'hbd) ?
                          reg826 : forvar842)) : $signed($unsigned(forvar826))) && ($signed(reg835) ^ forvar838)));
            end
          if ((($unsigned($unsigned($unsigned(wire823))) ?
                  $signed(forvar838) : reg841) ?
              reg826 : ((((~^wire821) != reg839[(1'h0):(1'h0)]) >= (~&(reg828 && reg832))) ?
                  "PO9odxOR" : reg830[(3'h4):(1'h1)])))
            begin
              reg850 <= forvar826;
              reg851 = wire822;
              reg852 = reg849;
              reg853 = wire824[(3'h4):(3'h4)];
              reg854 <= reg836[(4'ha):(4'h8)];
            end
          else
            begin
              reg850 = reg827;
              reg851 = wire824;
            end
        end
      if (forvar842[(2'h3):(1'h0)])
        begin
          for (forvar855 = (1'h0); (forvar855 < (1'h0)); forvar855 = (forvar855 + (1'h1)))
            begin
              reg856 <= (!reg844);
              reg857 <= {((&reg840[(2'h3):(2'h3)]) ?
                      reg841 : $unsigned(reg831[(2'h3):(2'h2)])),
                  (|(wire824 ?
                      (wire821[(3'h7):(3'h5)] ?
                          forvar838 : (reg853 * reg839)) : forvar826))};
              reg858 <= (reg827 ? forvar842 : forvar843[(4'he):(3'h5)]);
              reg859 = reg828;
              reg860 <= (($unsigned(((forvar832 * reg846) ^~ (forvar842 ?
                      reg844 : (8'hb0)))) ?
                  ((7'h44) ?
                      reg853 : ((reg858 && (8'ha4)) ?
                          (^~forvar827) : reg834[(1'h1):(1'h0)])) : $signed($unsigned($unsigned(reg841)))) ^ $unsigned({(8'h9d),
                  forvar835}));
            end
          if ({(reg859 ?
                  $unsigned($unsigned((!wire820))) : (forvar829 > $signed($signed((8'hb5))))),
              $signed(((&$unsigned(reg828)) ?
                  $signed({forvar826}) : reg829[(3'h4):(3'h4)]))})
            begin
              reg861 <= $signed($signed(($signed($unsigned(reg851)) > {$signed(wire824)})));
              reg862 = (forvar831[(4'h9):(4'h9)] << $signed(forvar829));
              reg863 = {reg858, {$signed(reg831), "U5FXta4OsJF"}};
              reg864 = reg863[(3'h6):(2'h2)];
              reg865 <= (~$unsigned((8'hbd)));
            end
          else
            begin
              reg861 <= $signed(reg862);
              reg862 <= ({(^((+forvar832) ? $unsigned(forvar842) : (|reg849))),
                  ($signed((!reg827)) & (^$unsigned(reg828)))} == $signed((+$signed($unsigned((8'hb9))))));
              reg863 <= forvar831[(3'h7):(2'h3)];
              reg864 <= $signed(wire822[(4'h9):(3'h5)]);
            end
          reg866 <= $unsigned(reg865);
        end
      else
        begin
          reg855 <= ($signed($unsigned(forvar826[(4'h9):(4'h9)])) ?
              reg845 : ({($signed((8'hbf)) ?
                      (~(8'hbc)) : (reg841 ? (7'h43) : reg841)),
                  {(reg829 ? (8'haf) : reg840), (reg848 * reg853)}} ^~ reg845));
        end
      for (forvar867 = (1'h0); (forvar867 < (1'h0)); forvar867 = (forvar867 + (1'h1)))
        begin
          reg868 = ($unsigned("fGrHBBfZzz5NFWSNo") == (reg832[(4'ha):(3'h7)] || $signed(reg856[(3'h6):(3'h5)])));
          for (forvar869 = (1'h0); (forvar869 < (1'h1)); forvar869 = (forvar869 + (1'h1)))
            begin
              reg870 = $unsigned("03");
            end
          reg871 <= $unsigned($unsigned($signed($unsigned($signed(forvar843)))));
          for (forvar872 = (1'h0); (forvar872 < (2'h3)); forvar872 = (forvar872 + (1'h1)))
            begin
              reg873 = (!reg865[(3'h4):(1'h0)]);
              reg874 = $signed((reg829[(3'h4):(2'h2)] ?
                  $unsigned(reg860) : (($unsigned(reg865) ^ forvar827[(1'h0):(1'h0)]) << wire820[(4'h8):(3'h6)])));
              reg875 = {$unsigned($signed($signed((forvar842 ~^ reg871)))),
                  "xYRZGLxwcUQZid"};
              reg876 <= (~^((-(forvar872 ?
                      {reg830, (8'hb8)} : $unsigned(reg853))) ?
                  (!((reg828 < reg831) ?
                      (reg851 ? forvar843 : reg829) : (wire825 ?
                          reg832 : reg850))) : forvar826));
              reg877 = (reg855 == forvar826[(1'h0):(1'h0)]);
            end
          reg878 <= ($signed({$signed($unsigned(reg857)),
              reg850}) || ((~^{$unsigned(forvar838), $signed(reg835)}) ?
              $signed(reg833) : reg848[(1'h0):(1'h0)]));
        end
      reg879 <= $signed((8'hbb));
    end
  assign wire880 = (~$signed(wire822));
  always
    @(posedge clk) begin
      for (forvar881 = (1'h0); (forvar881 < (2'h2)); forvar881 = (forvar881 + (1'h1)))
        begin
          reg882 <= "w3yUr3yfiNWPmW";
          if ((forvar832 ?
              $signed({((^wire821) ? $unsigned(reg845) : reg854[(3'h7):(3'h4)]),
                  {{reg850, reg837}, $unsigned(reg849)}}) : (!(|({reg882,
                  reg877} + $unsigned(reg862))))))
            begin
              reg883 = (|(~(&$unsigned(forvar869[(3'h5):(1'h0)]))));
              reg884 <= $signed((^reg844));
              reg885 <= {$unsigned($signed(wire825[(3'h5):(1'h1)]))};
              reg886 <= (-((reg863[(3'h6):(2'h3)] ?
                      $signed($unsigned((8'ha4))) : forvar832) ?
                  $unsigned(reg876[(5'h10):(4'hf)]) : (~^((~reg885) ?
                      ((8'ha4) >> reg862) : {reg847, (8'hb4)}))));
              reg887 <= reg886[(3'h5):(1'h1)];
            end
          else
            begin
              reg883 = ({forvar872[(1'h0):(1'h0)]} ?
                  reg887[(2'h3):(1'h1)] : (reg840 ~^ (((+forvar872) ?
                          (reg835 ? reg853 : reg874) : $unsigned(reg861)) ?
                      reg845[(3'h4):(1'h0)] : $signed($unsigned(reg878)))));
              reg884 <= $unsigned((reg855[(3'h4):(2'h2)] - ((reg873 ?
                  reg834 : "slT2") - ((forvar838 ?
                  reg870 : reg836) ^ reg840[(3'h5):(3'h5)]))));
              reg885 <= reg844;
              reg886 <= {reg874};
            end
        end
      reg888 <= (~&(~|(~|(|(-(7'h44))))));
    end
  assign wire889 = reg885[(3'h6):(2'h2)];
  assign wire890 = reg834[(4'h9):(3'h5)];
  assign wire891 = (~^$unsigned((((reg882 <<< wire819) ?
                           wire822[(3'h7):(1'h0)] : $signed(wire890)) ?
                       ("Br" <<< forvar842[(4'hc):(3'h4)]) : (^reg884[(1'h0):(1'h0)]))));
  assign wire892 = (reg840 != (forvar826[(3'h7):(3'h6)] ?
                       ((!(reg857 <<< (8'h9f))) ?
                           (forvar832 ?
                               {reg830,
                                   reg885} : (-reg851)) : ($unsigned((8'hba)) >= (reg862 >>> forvar827))) : reg870[(3'h4):(1'h1)]));
  assign wire893 = reg855[(1'h0):(1'h0)];
  assign wire894 = reg827[(3'h5):(3'h4)];
  assign wire895 = $unsigned(forvar829[(4'hc):(2'h3)]);
  assign wire896 = ({reg850[(5'h12):(4'hb)]} >>> {reg847,
                       $signed(($signed(wire894) ?
                           $signed(forvar843) : $unsigned(reg882)))});
  always
    @(posedge clk) begin
      if (($unsigned($unsigned($unsigned(forvar881[(4'ha):(1'h0)]))) ^~ reg828))
        begin
          for (forvar897 = (1'h0); (forvar897 < (2'h2)); forvar897 = (forvar897 + (1'h1)))
            begin
              reg898 <= reg884[(1'h1):(1'h0)];
              reg899 <= (reg887 + reg860);
              reg900 <= reg856[(4'h8):(2'h3)];
              reg901 <= $unsigned((~$signed((~^(^wire893)))));
            end
        end
      else
        begin
          for (forvar897 = (1'h0); (forvar897 < (1'h1)); forvar897 = (forvar897 + (1'h1)))
            begin
              reg898 <= (|((($unsigned(wire825) ?
                      $unsigned(reg849) : reg875[(2'h2):(2'h2)]) ?
                  ({reg840, reg871} ?
                      reg847 : {wire824}) : ((reg888 ^~ (8'ha7)) ~^ (forvar826 ?
                      reg862 : reg833))) > reg834));
              reg899 <= $signed(reg848[(1'h0):(1'h0)]);
              reg900 <= (~&$signed($signed(reg886[(4'hb):(3'h7)])));
              reg901 <= $signed($signed(reg882[(2'h2):(1'h1)]));
              reg902 = reg840[(4'hb):(2'h2)];
            end
          for (forvar903 = (1'h0); (forvar903 < (1'h1)); forvar903 = (forvar903 + (1'h1)))
            begin
              reg904 = (~$signed($signed($signed(reg857))));
              reg905 <= $unsigned({{(+$signed(forvar897))},
                  (forvar835 - $unsigned($signed(forvar855)))});
              reg906 <= ((($unsigned({forvar838,
                      reg859}) > ((~reg866) != (reg848 != reg850))) | (((forvar869 ?
                      reg886 : wire890) << $signed((8'ha1))) && (+{forvar843}))) ?
                  (reg833[(2'h3):(1'h1)] ?
                      $unsigned(((reg857 ? forvar872 : reg844) ?
                          (+reg834) : reg830)) : (~$signed(reg888))) : $signed((^~reg847[(3'h7):(1'h0)])));
            end
          reg907 = $unsigned(wire896);
          reg908 <= $unsigned($signed($unsigned((~^(8'hb9)))));
          for (forvar909 = (1'h0); (forvar909 < (1'h0)); forvar909 = (forvar909 + (1'h1)))
            begin
              reg910 = "Sh7coUZYBFxlkQSfPv";
              reg911 <= (8'haf);
            end
        end
      reg912 = ({reg904[(1'h1):(1'h1)]} < ((reg862[(4'h9):(2'h3)] <= ((-wire895) ?
              {reg849} : $signed(reg839))) ?
          (wire819[(4'h9):(3'h4)] >> reg827) : forvar826));
      reg913 = reg858[(4'ha):(3'h5)];
      reg914 = (reg913 << (-forvar838));
      if ($unsigned((8'ha4)))
        begin
          for (forvar915 = (1'h0); (forvar915 < (1'h1)); forvar915 = (forvar915 + (1'h1)))
            begin
              reg916 <= ($unsigned(((reg901 ?
                      (reg913 ?
                          forvar855 : forvar827) : (8'hb4)) | reg913[(3'h4):(1'h0)])) ?
                  wire822 : $unsigned($signed({(reg827 | reg904),
                      $signed((8'hb9))})));
              reg917 <= ($unsigned((8'had)) > $signed({((wire823 + forvar855) ?
                      $signed(reg837) : wire821[(4'h9):(1'h1)]),
                  (wire893 ? ((8'hb5) & reg908) : (~&wire824))}));
              reg918 <= (8'hb2);
            end
          reg919 <= $signed((&$signed($unsigned(reg837))));
          reg920 = {$signed((8'h9d))};
          reg921 = $unsigned(($signed($signed($signed(reg850))) + wire889));
          reg922 = $unsigned($unsigned(({reg905} != $signed((forvar832 ?
              forvar843 : wire891)))));
        end
      else
        begin
          for (forvar915 = (1'h0); (forvar915 < (3'h4)); forvar915 = (forvar915 + (1'h1)))
            begin
              reg916 = forvar855;
              reg917 <= $unsigned(($signed(reg863[(2'h3):(2'h2)]) ?
                  (reg866[(1'h1):(1'h0)] > {(reg887 < forvar897),
                      $unsigned(forvar842)}) : (reg855[(2'h2):(1'h0)] && reg914[(5'h12):(4'h9)])));
              reg918 <= $unsigned(reg870[(2'h2):(1'h0)]);
              reg919 = $unsigned(((+($signed(forvar831) ?
                  $signed(reg874) : (forvar903 ? reg849 : reg836))) || reg901));
            end
          if (({(({reg865} || reg911[(1'h1):(1'h1)]) >= reg879[(1'h1):(1'h0)])} != ($unsigned(reg913[(3'h6):(2'h2)]) | ((reg848[(1'h0):(1'h0)] != (reg849 ^ reg888)) > $unsigned($signed((8'hb3)))))))
            begin
              reg920 <= {reg841};
              reg921 <= $unsigned($signed((-($signed(reg873) ?
                  (forvar835 ? reg826 : reg849) : (reg863 ?
                      (7'h42) : forvar903)))));
            end
          else
            begin
              reg920 = "5dG7egD";
              reg921 = {$unsigned((8'haa)), (~forvar872[(1'h0):(1'h0)])};
            end
          for (forvar922 = (1'h0); (forvar922 < (3'h4)); forvar922 = (forvar922 + (1'h1)))
            begin
              reg923 <= reg873;
              reg924 <= (($unsigned($unsigned((reg841 ? reg899 : reg877))) ?
                      $unsigned($signed((reg826 ?
                          reg831 : reg901))) : (&{(wire880 ?
                              forvar835 : forvar827),
                          (^~reg875)})) ?
                  ({$unsigned((~&reg920))} + (!reg868[(4'he):(4'ha)])) : reg922[(4'hf):(3'h7)]);
              reg925 <= (reg900 ?
                  ("F0M0YUkq1VOQav" ?
                      {{$unsigned(forvar872)}} : $signed((~|$unsigned((8'hb7))))) : reg866);
              reg926 = $signed(((&reg849[(4'ha):(3'h4)]) == (forvar897[(1'h1):(1'h0)] ?
                  "9NNvG" : $signed((reg850 ^~ reg882)))));
              reg927 <= ((8'ha4) >> forvar872[(2'h2):(1'h1)]);
            end
          reg928 = (reg835[(3'h6):(1'h0)] ?
              "CCWFXU" : ((~&{forvar872[(1'h0):(1'h0)],
                      forvar867[(3'h7):(2'h2)]}) ?
                  $unsigned(($signed(reg847) ?
                      $signed(forvar832) : $unsigned(forvar832))) : $signed(($signed(reg913) ?
                      (&forvar881) : $signed(reg837)))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar929 = (1'h0); (forvar929 < (3'h4)); forvar929 = (forvar929 + (1'h1)))
        begin
          for (forvar930 = (1'h0); (forvar930 < (1'h1)); forvar930 = (forvar930 + (1'h1)))
            begin
              reg931 = (^(~|(forvar903 ? forvar827[(1'h1):(1'h0)] : reg888)));
              reg932 <= $signed({"4e0o1SgcAJovfeUvu",
                  (($signed(forvar842) > reg844[(4'h8):(1'h1)]) ?
                      ($unsigned(forvar909) >>> $unsigned(reg879)) : $signed((wire894 & forvar826)))});
              reg933 <= (("UrAmp6qE" ?
                  reg919[(3'h6):(3'h6)] : "hR9") + $signed(((|$unsigned((8'h9c))) < reg849[(3'h7):(1'h1)])));
              reg934 = {$signed($signed(reg873))};
            end
          reg935 <= $unsigned(reg846);
          for (forvar936 = (1'h0); (forvar936 < (1'h1)); forvar936 = (forvar936 + (1'h1)))
            begin
              reg937 <= (wire819 ?
                  reg838[(2'h3):(1'h1)] : $unsigned($unsigned(reg927[(3'h5):(2'h2)])));
              reg938 <= reg866;
            end
          for (forvar939 = (1'h0); (forvar939 < (3'h4)); forvar939 = (forvar939 + (1'h1)))
            begin
              reg940 <= forvar903[(4'h9):(3'h6)];
              reg941 = (reg898 ?
                  forvar832[(3'h4):(2'h3)] : {(reg866 < {forvar936}),
                      {wire880[(3'h6):(3'h4)], reg868}});
              reg942 <= (wire819[(4'ha):(4'ha)] >> (($signed(forvar832[(2'h2):(2'h2)]) ?
                  {$signed(reg845),
                      (reg844 ? wire891 : wire892)} : $signed(((8'ha7) ?
                      (8'hbd) : reg826))) && (({reg926, (8'hbf)} ?
                  {forvar929} : $signed(reg866)) || $signed($unsigned((8'hb1))))));
            end
        end
      for (forvar943 = (1'h0); (forvar943 < (1'h0)); forvar943 = (forvar943 + (1'h1)))
        begin
          reg944 <= ($unsigned({({(8'hb3)} ?
                  reg834[(4'hb):(3'h6)] : (^(7'h40)))}) > wire891);
          if ((reg907 ^~ $unsigned($signed($signed((&reg838))))))
            begin
              reg945 <= $unsigned((^~(reg868 - {wire819[(3'h7):(1'h1)],
                  wire893[(4'hb):(3'h7)]})));
              reg946 <= forvar939[(3'h7):(1'h0)];
              reg947 <= {reg934[(2'h2):(2'h2)],
                  (($unsigned($signed(reg831)) ?
                          $signed((!reg925)) : ((^~reg857) | wire819)) ?
                      $unsigned(((wire822 >>> (8'haf)) - wire894[(4'h8):(2'h2)])) : "mPcJquCab8RCMVSl")};
            end
          else
            begin
              reg945 <= wire891;
              reg946 <= $signed((($unsigned((~reg828)) ?
                      $unsigned((+wire824)) : ($signed(reg877) ?
                          (reg942 > reg926) : reg912[(5'h15):(4'hf)])) ?
                  (8'hb0) : (&$signed($signed(reg877)))));
              reg947 = $unsigned(forvar922);
            end
          for (forvar948 = (1'h0); (forvar948 < (1'h0)); forvar948 = (forvar948 + (1'h1)))
            begin
              reg949 <= (8'ha5);
              reg950 = reg901[(3'h4):(3'h4)];
            end
        end
      for (forvar951 = (1'h0); (forvar951 < (1'h1)); forvar951 = (forvar951 + (1'h1)))
        begin
          for (forvar952 = (1'h0); (forvar952 < (1'h0)); forvar952 = (forvar952 + (1'h1)))
            begin
              reg953 <= ({(~reg902[(3'h5):(1'h1)]),
                  {((reg840 ? reg839 : reg906) > reg827),
                      ((~reg865) ?
                          (reg833 ~^ reg919) : {wire892,
                              reg856})}} ~^ ("uRn" ~^ reg854));
              reg954 <= {$unsigned(forvar922[(3'h5):(3'h4)])};
              reg955 <= ((8'ha0) ?
                  {reg868,
                      (reg826 ?
                          $unsigned($unsigned(reg849)) : $unsigned((reg888 ?
                              reg838 : reg848)))} : (reg829 ?
                      ((&(wire892 ? (8'hb8) : reg846)) ?
                          reg928[(4'hc):(3'h6)] : $signed({reg899,
                              (7'h40)})) : $signed(reg913)));
            end
          reg956 = forvar881;
          for (forvar957 = (1'h0); (forvar957 < (1'h0)); forvar957 = (forvar957 + (1'h1)))
            begin
              reg958 <= reg953[(2'h3):(2'h3)];
              reg959 <= reg908;
              reg960 <= (-(($unsigned($signed(forvar838)) ~^ ($signed(reg884) == (reg844 << reg956))) ?
                  $signed($signed((reg918 + forvar909))) : ((^{reg833}) & reg912[(4'h8):(3'h5)])));
              reg961 = reg850;
            end
          for (forvar962 = (1'h0); (forvar962 < (1'h1)); forvar962 = (forvar962 + (1'h1)))
            begin
              reg963 = (((|reg910[(3'h5):(2'h2)]) ?
                      reg961[(5'h13):(5'h12)] : (&(-$unsigned((8'haa))))) ?
                  reg904 : $unsigned((reg859 ? reg942 : (^~reg833))));
            end
          for (forvar964 = (1'h0); (forvar964 < (1'h0)); forvar964 = (forvar964 + (1'h1)))
            begin
              reg965 = forvar869;
            end
        end
      reg966 = reg956[(5'h11):(1'h1)];
      for (forvar967 = (1'h0); (forvar967 < (1'h1)); forvar967 = (forvar967 + (1'h1)))
        begin
          if (($unsigned({reg871}) ?
              $signed((reg850 ?
                  {$unsigned(reg926)} : ($unsigned(reg885) * $unsigned((8'ha0))))) : ((~|reg906) ?
                  $signed((+reg935)) : (^~$signed(((8'hb8) && forvar838))))))
            begin
              reg968 = ($unsigned($signed(reg850[(3'h7):(3'h4)])) ?
                  {((reg931[(1'h1):(1'h1)] ?
                          (reg938 ? reg888 : reg826) : {wire890,
                              reg884}) & (7'h44)),
                      (8'hbf)} : (~($unsigned($signed(wire894)) ?
                      reg845[(2'h2):(2'h2)] : (^~$signed(reg888)))));
              reg969 <= $unsigned($signed($unsigned((wire889[(1'h1):(1'h1)] ?
                  reg942 : $unsigned(reg966)))));
              reg970 <= (^~reg863[(4'hb):(4'h8)]);
              reg971 = $unsigned($signed(reg826[(4'hc):(4'h8)]));
              reg972 <= {(|$unsigned((+reg898)))};
            end
          else
            begin
              reg968 <= forvar855;
              reg969 <= ((^~forvar881) ?
                  (reg950 ?
                      $unsigned({(~^reg956),
                          $unsigned(reg912)}) : (~^reg944[(4'hf):(4'h9)])) : (|$signed(reg933)));
              reg970 <= {(($signed($signed(reg840)) && ((reg838 ?
                          reg844 : reg856) >= (reg925 & reg971))) ?
                      ($signed("4D3") ?
                          (^~reg924[(2'h2):(2'h2)]) : ((reg960 ?
                              reg827 : reg938) ^ ((8'hb6) + reg935))) : (forvar827 ?
                          reg878 : $unsigned($signed(wire892)))),
                  (-{(~$signed(reg836))})};
              reg971 <= {$unsigned({reg947[(1'h0):(1'h0)], reg847})};
            end
          for (forvar973 = (1'h0); (forvar973 < (2'h2)); forvar973 = (forvar973 + (1'h1)))
            begin
              reg974 <= (!$unsigned(((reg947 ? $unsigned(reg868) : (8'h9c)) ?
                  ($unsigned(reg844) ?
                      (wire896 ?
                          reg934 : (8'h9e)) : (forvar952 ^ forvar842)) : ($unsigned(reg906) * (reg931 <<< reg907)))));
            end
          reg975 = reg838[(1'h0):(1'h0)];
        end
    end
  assign wire976 = reg862;
  always
    @(posedge clk) begin
      reg977 = (reg904 ?
          (&$unsigned(forvar826[(3'h7):(1'h0)])) : "Al181XqPHQhaiv7AsEU0");
      for (forvar978 = (1'h0); (forvar978 < (2'h3)); forvar978 = (forvar978 + (1'h1)))
        begin
          for (forvar979 = (1'h0); (forvar979 < (1'h1)); forvar979 = (forvar979 + (1'h1)))
            begin
              reg980 <= ($unsigned($unsigned((forvar978[(5'h10):(3'h4)] ?
                  (reg913 ?
                      forvar948 : wire893) : (8'hb2)))) && ($unsigned((8'h9c)) <<< $signed({reg839})));
              reg981 <= reg914[(4'hb):(1'h1)];
              reg982 <= reg931[(2'h2):(1'h1)];
              reg983 <= reg898;
              reg984 <= $signed($unsigned($signed($signed($unsigned(reg956)))));
            end
          reg985 <= (reg839[(5'h10):(4'hf)] << ({{forvar832[(2'h2):(2'h2)]}} - reg969[(3'h6):(2'h2)]));
          for (forvar986 = (1'h0); (forvar986 < (2'h2)); forvar986 = (forvar986 + (1'h1)))
            begin
              reg987 <= $unsigned({$signed($unsigned((reg877 ^~ (8'hae))))});
              reg988 <= ($unsigned((wire976 ?
                  reg969 : ((reg908 >>> forvar903) & {forvar826,
                      forvar936}))) || (((|(reg851 ?
                      reg983 : reg882)) || ($unsigned(reg840) >> (+forvar957))) ?
                  {$unsigned((reg850 + reg932))} : reg922));
            end
          reg989 <= forvar855;
        end
      for (forvar990 = (1'h0); (forvar990 < (2'h3)); forvar990 = (forvar990 + (1'h1)))
        begin
          for (forvar991 = (1'h0); (forvar991 < (1'h1)); forvar991 = (forvar991 + (1'h1)))
            begin
              reg992 <= {forvar948};
            end
          for (forvar993 = (1'h0); (forvar993 < (2'h2)); forvar993 = (forvar993 + (1'h1)))
            begin
              reg994 <= wire821;
              reg995 <= (($unsigned($signed(reg983)) <<< reg912) ?
                  (^(|($unsigned(reg871) ?
                      $signed(reg859) : ((8'hbe) ?
                          reg845 : (8'ha2))))) : reg923[(2'h2):(1'h0)]);
              reg996 = reg834;
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module644
#( parameter param743 = {((({(8'hb9)} << ((8'hb9) ? (8'hba) : (8'ha9))) ? {((7'h44) ? (8'hab) : (8'ha4))} : (((8'hb6) >> (7'h40)) ? (^~(8'hb8)) : ((8'ha3) < (8'hbd)))) && (|(((7'h41) ? (8'haf) : (7'h43)) ? {(8'h9f), (7'h44)} : (7'h42)))), {(&(((8'hbe) ? (8'h9e) : (8'h9e)) != ((7'h43) > (8'ha7)))), (!(-((7'h40) >> (8'h9e))))}}
, parameter param744 = (((-param743) ? (&(~&{param743})) : param743) >> {(8'had)}) )
(y, clk, wire648, wire647, wire646, wire645);
  output wire [(32'h451):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire648;
  input wire [(5'h10):(1'h0)] wire647;
  input wire [(5'h11):(1'h0)] wire646;
  input wire [(4'hd):(1'h0)] wire645;
  wire [(4'hf):(1'h0)] wire742;
  reg [(5'h14):(1'h0)] reg741 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg740 = (1'h0);
  reg [(4'hf):(1'h0)] reg739 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar738 = (1'h0);
  reg [(5'h13):(1'h0)] reg737 = (1'h0);
  reg [(3'h5):(1'h0)] reg736 = (1'h0);
  wire [(3'h5):(1'h0)] wire735;
  wire [(4'hd):(1'h0)] wire734;
  wire [(5'h12):(1'h0)] wire733;
  reg [(5'h12):(1'h0)] reg732 = (1'h0);
  reg [(5'h12):(1'h0)] reg731 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg730 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar729 = (1'h0);
  reg [(5'h15):(1'h0)] reg728 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg727 = (1'h0);
  reg [(4'ha):(1'h0)] reg726 = (1'h0);
  reg [(3'h4):(1'h0)] reg725 = (1'h0);
  reg [(4'hd):(1'h0)] reg724 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar723 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar722 = (1'h0);
  reg [(2'h3):(1'h0)] reg721 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg720 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar719 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg718 = (1'h0);
  reg [(4'ha):(1'h0)] reg717 = (1'h0);
  reg [(5'h12):(1'h0)] reg716 = (1'h0);
  reg [(2'h2):(1'h0)] reg715 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar714 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg713 = (1'h0);
  reg [(2'h2):(1'h0)] reg712 = (1'h0);
  reg [(4'hf):(1'h0)] reg711 = (1'h0);
  reg [(4'h9):(1'h0)] reg710 = (1'h0);
  reg [(5'h10):(1'h0)] reg709 = (1'h0);
  reg [(4'h8):(1'h0)] forvar708 = (1'h0);
  reg [(4'hf):(1'h0)] reg707 = (1'h0);
  reg signed [(4'he):(1'h0)] reg706 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg705 = (1'h0);
  reg [(2'h3):(1'h0)] reg704 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar703 = (1'h0);
  reg [(5'h10):(1'h0)] reg702 = (1'h0);
  reg [(5'h13):(1'h0)] reg701 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg700 = (1'h0);
  reg [(4'hd):(1'h0)] reg699 = (1'h0);
  reg [(5'h14):(1'h0)] reg698 = (1'h0);
  reg [(5'h10):(1'h0)] forvar697 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar696 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg695 = (1'h0);
  reg [(4'hd):(1'h0)] reg694 = (1'h0);
  reg [(5'h13):(1'h0)] reg693 = (1'h0);
  reg [(5'h11):(1'h0)] reg692 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg691 = (1'h0);
  reg [(3'h5):(1'h0)] reg690 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar689 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar688 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg687 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg686 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg685 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg684 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg683 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg682 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar681 = (1'h0);
  reg [(4'hf):(1'h0)] reg680 = (1'h0);
  reg [(4'h9):(1'h0)] forvar679 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar678 = (1'h0);
  wire signed [(3'h6):(1'h0)] wire677;
  reg signed [(4'hf):(1'h0)] reg676 = (1'h0);
  reg [(4'ha):(1'h0)] forvar669 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg668 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg675 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg674 = (1'h0);
  reg [(2'h3):(1'h0)] reg673 = (1'h0);
  reg [(4'hb):(1'h0)] reg672 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg671 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg670 = (1'h0);
  reg [(4'hc):(1'h0)] reg669 = (1'h0);
  reg [(5'h11):(1'h0)] forvar668 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg667 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg666 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg664 = (1'h0);
  reg [(5'h10):(1'h0)] reg663 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg662 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg661 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar660 = (1'h0);
  reg [(4'ha):(1'h0)] forvar659 = (1'h0);
  reg [(5'h11):(1'h0)] reg658 = (1'h0);
  reg [(4'h9):(1'h0)] reg657 = (1'h0);
  reg [(4'h9):(1'h0)] forvar656 = (1'h0);
  wire signed [(3'h5):(1'h0)] wire655;
  wire signed [(5'h14):(1'h0)] wire654;
  wire signed [(3'h7):(1'h0)] wire653;
  wire [(4'hd):(1'h0)] wire652;
  reg signed [(3'h7):(1'h0)] reg651 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire650;
  wire signed [(5'h11):(1'h0)] wire649;
  assign y = {wire742,
                 reg741,
                 reg740,
                 reg739,
                 forvar738,
                 reg737,
                 reg736,
                 wire735,
                 wire734,
                 wire733,
                 reg732,
                 reg731,
                 reg730,
                 forvar729,
                 reg728,
                 reg727,
                 reg726,
                 reg725,
                 reg724,
                 forvar723,
                 forvar722,
                 reg721,
                 reg720,
                 forvar719,
                 reg718,
                 reg717,
                 reg716,
                 reg715,
                 forvar714,
                 reg713,
                 reg712,
                 reg711,
                 reg710,
                 reg709,
                 forvar708,
                 reg707,
                 reg706,
                 reg705,
                 reg704,
                 forvar703,
                 reg702,
                 reg701,
                 reg700,
                 reg699,
                 reg698,
                 forvar697,
                 forvar696,
                 reg695,
                 reg694,
                 reg693,
                 reg692,
                 reg691,
                 reg690,
                 forvar689,
                 forvar688,
                 reg687,
                 reg686,
                 reg685,
                 reg684,
                 reg683,
                 reg682,
                 forvar681,
                 reg680,
                 forvar679,
                 forvar678,
                 wire677,
                 reg676,
                 forvar669,
                 reg668,
                 reg675,
                 reg674,
                 reg673,
                 reg672,
                 reg671,
                 reg670,
                 reg669,
                 forvar668,
                 reg667,
                 reg666,
                 reg665,
                 reg664,
                 reg663,
                 reg662,
                 reg661,
                 forvar660,
                 forvar659,
                 reg658,
                 reg657,
                 forvar656,
                 wire655,
                 wire654,
                 wire653,
                 wire652,
                 reg651,
                 wire650,
                 wire649,
                 (1'h0)};
  assign wire649 = $unsigned(((~^($unsigned(wire647) && ((8'h9f) ?
                           wire648 : wire645))) ?
                       {($signed(wire647) ? wire646 : {wire645}),
                           (+(+(7'h40)))} : wire645[(4'hd):(3'h6)]));
  assign wire650 = $unsigned(wire648);
  always
    @(posedge clk) begin
      reg651 <= wire645;
    end
  assign wire652 = $signed((8'ha3));
  assign wire653 = ($signed($signed(($unsigned(wire648) ?
                       (wire646 ?
                           wire645 : wire645) : wire652[(3'h6):(2'h2)]))) >> (~&(wire646 ?
                       ((wire647 >> wire645) > (wire648 || wire652)) : $unsigned({wire646,
                           (8'hbe)}))));
  assign wire654 = wire649;
  assign wire655 = (-$signed({wire646, $signed($unsigned(wire653))}));
  always
    @(posedge clk) begin
      for (forvar656 = (1'h0); (forvar656 < (1'h0)); forvar656 = (forvar656 + (1'h1)))
        begin
          reg657 <= $signed(wire649[(4'ha):(4'h9)]);
          reg658 <= (^"bNmbcmHtC");
        end
    end
  always
    @(posedge clk) begin
      for (forvar659 = (1'h0); (forvar659 < (2'h2)); forvar659 = (forvar659 + (1'h1)))
        begin
          for (forvar660 = (1'h0); (forvar660 < (2'h2)); forvar660 = (forvar660 + (1'h1)))
            begin
              reg661 = {$signed((~(forvar660[(2'h3):(1'h0)] >>> ((8'hae) < wire647)))),
                  (($unsigned(wire655) ?
                      "F1Y5mZ5IwmAeZ8" : (8'ha2)) << (7'h42))};
              reg662 <= ((+(^~$unsigned((reg661 << wire648)))) <<< $signed(((8'h9f) ?
                  {wire654[(5'h14):(4'hf)]} : (^(+wire648)))));
              reg663 = ((~wire655[(1'h0):(1'h0)]) * {reg658});
            end
          reg664 = {"eIPoapb", $unsigned(reg661)};
          reg665 = (+$signed(wire648));
          reg666 <= ($signed(((reg663[(4'h9):(1'h0)] * forvar660) ?
                  ($unsigned(wire654) << $unsigned(forvar660)) : $signed((-wire653)))) ?
              reg663[(3'h7):(1'h1)] : ((!$signed((~^wire653))) ?
                  reg661 : $signed(($signed((8'hb5)) << $signed(wire653)))));
        end
      reg667 <= (wire647[(3'h4):(1'h1)] ?
          ($unsigned(($signed(wire645) ?
              (reg657 + forvar656) : $unsigned(wire647))) && $unsigned($unsigned((reg658 ?
              wire652 : reg658)))) : $signed((({wire650} * reg661) ?
              {wire646} : $unsigned((-forvar656)))));
      if (wire649[(4'h8):(3'h7)])
        begin
          for (forvar668 = (1'h0); (forvar668 < (1'h0)); forvar668 = (forvar668 + (1'h1)))
            begin
              reg669 = wire647[(4'hd):(4'h8)];
              reg670 = ((+$signed($signed((reg667 ~^ (8'hb1))))) ?
                  reg665 : forvar659);
            end
          if (wire647[(1'h1):(1'h0)])
            begin
              reg671 <= (8'ha1);
              reg672 = reg662;
            end
          else
            begin
              reg671 <= (wire653[(3'h4):(1'h0)] ?
                  $unsigned({(reg658 & (reg661 ?
                          wire652 : reg665))}) : ((wire647[(4'hb):(1'h1)] ?
                          wire655[(2'h2):(1'h0)] : (~$unsigned(reg651))) ?
                      (reg664[(3'h4):(2'h2)] ?
                          (&wire646[(4'hc):(4'h9)]) : (-reg662[(2'h2):(1'h1)])) : ($signed($unsigned((8'ha5))) == $signed((forvar656 ?
                          wire653 : reg665)))));
              reg672 <= (^$unsigned($signed($unsigned($signed(reg662)))));
              reg673 <= $unsigned(((reg665 + (~&(wire646 >> reg669))) > wire648));
              reg674 = wire649[(4'he):(3'h5)];
              reg675 <= wire647[(3'h5):(1'h1)];
            end
        end
      else
        begin
          reg668 <= $signed($unsigned({$signed($unsigned(wire648)), (8'hb3)}));
          for (forvar669 = (1'h0); (forvar669 < (2'h2)); forvar669 = (forvar669 + (1'h1)))
            begin
              reg670 = wire645;
              reg671 <= ($signed(wire654[(4'ha):(2'h3)]) ?
                  reg673[(1'h0):(1'h0)] : $unsigned(reg672));
              reg672 = $unsigned((!(reg666[(2'h2):(1'h0)] | {(reg664 ?
                      reg672 : wire650),
                  reg662})));
              reg673 = $signed((+$signed($unsigned((~&forvar659)))));
            end
        end
      reg676 <= (reg667[(2'h2):(1'h1)] == ($unsigned($unsigned(forvar656[(3'h5):(2'h2)])) ?
          (((8'hbd) <<< (8'ha1)) > (8'hbf)) : reg664));
    end
  assign wire677 = (wire655 ?
                       (!reg675) : $signed(($signed((reg657 || reg651)) ?
                           {(reg669 ?
                                   reg658 : forvar669)} : $signed((8'ha4)))));
  always
    @(posedge clk) begin
      for (forvar678 = (1'h0); (forvar678 < (1'h1)); forvar678 = (forvar678 + (1'h1)))
        begin
          for (forvar679 = (1'h0); (forvar679 < (1'h1)); forvar679 = (forvar679 + (1'h1)))
            begin
              reg680 = $signed((+($signed("sX8") ^~ ($unsigned(reg658) ?
                  ((8'hae) ? forvar656 : (8'h9e)) : (^~forvar660)))));
            end
          for (forvar681 = (1'h0); (forvar681 < (2'h3)); forvar681 = (forvar681 + (1'h1)))
            begin
              reg682 <= ($signed((|(!(reg672 - forvar681)))) ?
                  ({$signed(forvar678), $signed((reg661 ? reg680 : wire652))} ?
                      {"OWSG9b5NQY9qU4E"} : (8'hb8)) : (((&(wire647 ?
                          reg669 : wire677)) == reg667) ?
                      $unsigned($unsigned({(8'h9e), wire655})) : wire646));
              reg683 <= "lA03lQz91l3JkF9N";
            end
          reg684 = forvar660;
          reg685 = reg668[(1'h0):(1'h0)];
          if ("qXZu")
            begin
              reg686 <= forvar679[(3'h5):(1'h1)];
              reg687 = reg685[(4'h8):(3'h6)];
            end
          else
            begin
              reg686 <= $unsigned((8'hbb));
              reg687 <= $signed($unsigned(wire649));
            end
        end
      for (forvar688 = (1'h0); (forvar688 < (2'h2)); forvar688 = (forvar688 + (1'h1)))
        begin
          for (forvar689 = (1'h0); (forvar689 < (2'h2)); forvar689 = (forvar689 + (1'h1)))
            begin
              reg690 = forvar668[(4'hd):(4'h9)];
              reg691 <= (~&("qbXcixW" ? reg669 : "cr8S"));
              reg692 <= $signed(((forvar689 ?
                  ({wire649} ?
                      (^~reg663) : $unsigned(reg675)) : {((8'h9c) >= (8'had)),
                      $signed(wire645)}) || (reg690[(2'h3):(2'h3)] ?
                  $unsigned((8'hb9)) : forvar679)));
            end
          reg693 <= {reg674[(3'h7):(3'h4)]};
          reg694 <= $unsigned(($signed(forvar689[(3'h7):(3'h5)]) ?
              $unsigned(((|wire646) | reg691[(2'h2):(2'h2)])) : $unsigned(($unsigned((8'ha4)) <= $signed(forvar688)))));
          reg695 = $unsigned(forvar660[(1'h1):(1'h1)]);
        end
      for (forvar696 = (1'h0); (forvar696 < (3'h4)); forvar696 = (forvar696 + (1'h1)))
        begin
          for (forvar697 = (1'h0); (forvar697 < (2'h2)); forvar697 = (forvar697 + (1'h1)))
            begin
              reg698 <= $signed($unsigned((-forvar681)));
              reg699 = $signed($signed((reg668[(3'h4):(2'h3)] > wire655)));
              reg700 <= reg698;
              reg701 <= $unsigned((($signed($signed(reg690)) ?
                      reg671 : ("BtVbcCtao" >> $signed((7'h43)))) ?
                  $signed((wire649[(4'hb):(3'h7)] ?
                      (~&(8'hb4)) : (reg666 & forvar696))) : ((reg662 <= {(8'ha1)}) >>> reg668[(3'h4):(1'h1)])));
              reg702 = ($signed(reg670) & forvar660);
            end
          for (forvar703 = (1'h0); (forvar703 < (2'h3)); forvar703 = (forvar703 + (1'h1)))
            begin
              reg704 = (-{"xB", {$unsigned(((8'ha8) ? wire654 : forvar660))}});
              reg705 = $unsigned($signed((8'h9e)));
              reg706 <= {$unsigned(($unsigned($unsigned(reg698)) >> reg682))};
            end
          reg707 <= (-$unsigned(reg671[(4'hf):(4'hd)]));
        end
      for (forvar708 = (1'h0); (forvar708 < (2'h2)); forvar708 = (forvar708 + (1'h1)))
        begin
          if ($signed((|{$unsigned($signed(forvar659))})))
            begin
              reg709 <= reg668;
            end
          else
            begin
              reg709 <= $signed(reg694);
              reg710 = {reg700[(2'h2):(1'h0)]};
              reg711 = (wire652[(3'h7):(2'h2)] ~^ (7'h40));
              reg712 <= {wire648[(2'h2):(1'h1)]};
              reg713 = ((^(~|$unsigned((~reg707)))) ?
                  $unsigned((!reg698[(2'h2):(1'h0)])) : reg662[(4'h9):(3'h4)]);
            end
          for (forvar714 = (1'h0); (forvar714 < (2'h3)); forvar714 = (forvar714 + (1'h1)))
            begin
              reg715 <= ($signed(((~&reg686[(2'h2):(1'h0)]) ?
                  {(forvar678 & wire653)} : $signed($unsigned(forvar681)))) >> ((reg692[(5'h10):(3'h4)] ?
                  reg682[(4'hb):(4'h9)] : ((reg693 * (7'h43)) ?
                      "G6ndNAllayTbkeMKs" : $signed(reg713))) != $unsigned(reg666)));
              reg716 = $signed((+{$unsigned(reg705[(3'h4):(2'h3)])}));
              reg717 <= $unsigned(reg707);
              reg718 <= (&forvar697[(1'h1):(1'h0)]);
            end
          for (forvar719 = (1'h0); (forvar719 < (3'h4)); forvar719 = (forvar719 + (1'h1)))
            begin
              reg720 <= {$signed(wire655[(3'h5):(3'h4)]), wire654};
            end
          reg721 <= wire677;
        end
      for (forvar722 = (1'h0); (forvar722 < (3'h4)); forvar722 = (forvar722 + (1'h1)))
        begin
          for (forvar723 = (1'h0); (forvar723 < (3'h4)); forvar723 = (forvar723 + (1'h1)))
            begin
              reg724 = wire645[(4'h9):(3'h6)];
              reg725 = forvar689;
              reg726 <= $signed((~&({forvar678, {wire654, reg716}} ?
                  (~{wire649}) : ("l" != (reg691 ^ forvar659)))));
            end
          reg727 = (((($unsigned(reg725) != reg701[(5'h13):(4'hd)]) ?
                  wire655 : {reg692}) ?
              (-$unsigned(reg706)) : (8'ha4)) | (((^~(^reg726)) ?
                  ($unsigned((8'had)) - reg682) : $unsigned({(8'ha3)})) ?
              $unsigned($signed({reg662})) : $unsigned((~&(8'hac)))));
          reg728 <= reg727[(2'h2):(2'h2)];
          for (forvar729 = (1'h0); (forvar729 < (1'h0)); forvar729 = (forvar729 + (1'h1)))
            begin
              reg730 = ((($unsigned((reg705 ?
                  forvar722 : reg668)) ~^ $unsigned((&reg665))) != forvar708[(3'h7):(1'h1)]) > {({((8'ha0) >> reg727),
                          forvar729} ?
                      (reg728 ?
                          reg658 : $unsigned((8'hac))) : {(forvar714 + forvar679),
                          forvar669})});
              reg731 <= (reg727 ?
                  reg657 : $unsigned($signed($unsigned((|reg666)))));
            end
          reg732 <= (reg720 || {reg692,
              (((forvar656 ? wire646 : forvar696) ?
                  (reg658 ? reg666 : wire652) : $signed(reg713)) > "n8ort")});
        end
    end
  assign wire733 = ($unsigned(((+$signed(reg699)) ?
                       ($signed(reg721) ?
                           forvar696[(3'h5):(1'h1)] : (reg712 >> (7'h43))) : forvar659)) ^ $unsigned((8'hbc)));
  assign wire734 = $unsigned((forvar703[(1'h0):(1'h0)] ?
                       {($signed(forvar696) > wire649),
                           reg685[(3'h5):(2'h3)]} : $unsigned(reg716[(5'h12):(5'h12)])));
  assign wire735 = reg686;
  always
    @(posedge clk) begin
      reg736 = (((reg676[(4'hf):(2'h3)] ?
          {$signed(wire733)} : $unsigned((|wire649))) > (~&reg695)) << forvar696[(3'h4):(3'h4)]);
      reg737 <= reg665[(3'h5):(3'h5)];
      for (forvar738 = (1'h0); (forvar738 < (3'h4)); forvar738 = (forvar738 + (1'h1)))
        begin
          if ({forvar719, $unsigned($unsigned("uphH2AWs5tlZYi"))})
            begin
              reg739 <= reg706;
              reg740 <= $signed((forvar660[(3'h4):(1'h1)] ?
                  reg670 : ($signed((~(8'h9f))) < ("5mw0TQ" == reg685))));
            end
          else
            begin
              reg739 <= forvar738[(1'h1):(1'h0)];
              reg740 <= ("" ?
                  ($signed($signed(wire734)) < reg713[(3'h5):(1'h1)]) : forvar688);
              reg741 = ((~^(reg686[(5'h12):(5'h10)] > (7'h41))) >>> wire649[(5'h11):(4'hd)]);
            end
        end
    end
  assign wire742 = (wire733 && (reg718 || forvar668[(3'h4):(2'h2)]));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module510
#( parameter param640 = ((~|{(!((8'h9c) ^~ (8'ha3))), (8'h9e)}) ? ((^{{(8'ha5)}}) ? ((~&(~|(8'ha1))) ? ({(8'ha3), (8'had)} < ((8'hb6) ? (8'hae) : (8'h9d))) : {(&(8'hb5))}) : (|(~&((8'haf) << (8'h9f))))) : (-{(~{(8'hb3)})}))
, parameter param641 = param640 )
(y, clk, wire515, wire514, wire513, wire512, wire511);
  output wire [(32'h5c2):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire515;
  input wire [(3'h7):(1'h0)] wire514;
  input wire [(3'h6):(1'h0)] wire513;
  input wire [(3'h6):(1'h0)] wire512;
  input wire [(3'h7):(1'h0)] wire511;
  wire [(4'h8):(1'h0)] wire639;
  wire signed [(3'h6):(1'h0)] wire638;
  wire [(5'h13):(1'h0)] wire637;
  wire signed [(4'h9):(1'h0)] wire636;
  wire signed [(3'h5):(1'h0)] wire635;
  wire signed [(4'hb):(1'h0)] wire634;
  wire signed [(2'h2):(1'h0)] wire633;
  wire signed [(5'h11):(1'h0)] wire632;
  wire signed [(2'h3):(1'h0)] wire631;
  reg [(5'h12):(1'h0)] reg630 = (1'h0);
  reg [(4'hf):(1'h0)] reg629 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg628 = (1'h0);
  reg [(3'h6):(1'h0)] forvar627 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg626 = (1'h0);
  reg [(2'h2):(1'h0)] reg625 = (1'h0);
  reg [(5'h14):(1'h0)] reg624 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg623 = (1'h0);
  reg [(5'h12):(1'h0)] reg622 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg621 = (1'h0);
  reg [(3'h6):(1'h0)] reg620 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar619 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar618 = (1'h0);
  reg [(3'h4):(1'h0)] reg614 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg617 = (1'h0);
  reg [(4'ha):(1'h0)] reg616 = (1'h0);
  reg [(4'hc):(1'h0)] reg615 = (1'h0);
  reg [(5'h15):(1'h0)] forvar614 = (1'h0);
  reg [(5'h14):(1'h0)] reg613 = (1'h0);
  reg [(5'h11):(1'h0)] reg612 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar611 = (1'h0);
  reg [(5'h10):(1'h0)] reg610 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar609 = (1'h0);
  reg [(4'ha):(1'h0)] reg608 = (1'h0);
  reg [(5'h11):(1'h0)] reg607 = (1'h0);
  wire signed [(4'h9):(1'h0)] wire606;
  wire [(5'h10):(1'h0)] wire605;
  reg [(3'h5):(1'h0)] reg604 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg603 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg602 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg601 = (1'h0);
  reg [(5'h13):(1'h0)] reg600 = (1'h0);
  reg [(4'hf):(1'h0)] forvar595 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar591 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg599 = (1'h0);
  reg [(2'h3):(1'h0)] reg598 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg597 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg596 = (1'h0);
  reg [(4'ha):(1'h0)] reg595 = (1'h0);
  reg [(2'h2):(1'h0)] reg594 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg593 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg592 = (1'h0);
  reg [(3'h5):(1'h0)] reg591 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg590 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg589 = (1'h0);
  reg [(5'h12):(1'h0)] reg588 = (1'h0);
  reg [(4'hb):(1'h0)] reg587 = (1'h0);
  reg [(3'h7):(1'h0)] forvar586 = (1'h0);
  reg [(2'h3):(1'h0)] reg585 = (1'h0);
  reg [(5'h14):(1'h0)] reg584 = (1'h0);
  reg [(5'h10):(1'h0)] reg583 = (1'h0);
  reg [(5'h14):(1'h0)] reg582 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg581 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg580 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar579 = (1'h0);
  wire signed [(3'h7):(1'h0)] wire578;
  wire [(2'h2):(1'h0)] wire577;
  reg signed [(5'h10):(1'h0)] forvar569 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg576 = (1'h0);
  reg [(5'h12):(1'h0)] reg575 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg574 = (1'h0);
  reg [(5'h10):(1'h0)] reg573 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar572 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg571 = (1'h0);
  reg signed [(4'he):(1'h0)] reg570 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg569 = (1'h0);
  reg [(4'hf):(1'h0)] reg568 = (1'h0);
  reg [(3'h5):(1'h0)] reg567 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg566 = (1'h0);
  reg [(5'h15):(1'h0)] forvar565 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg563 = (1'h0);
  reg [(3'h4):(1'h0)] reg562 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar561 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg560 = (1'h0);
  reg signed [(4'he):(1'h0)] reg559 = (1'h0);
  reg [(5'h12):(1'h0)] reg558 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire557;
  reg [(5'h14):(1'h0)] reg556 = (1'h0);
  reg [(4'hb):(1'h0)] reg555 = (1'h0);
  reg [(3'h6):(1'h0)] reg554 = (1'h0);
  reg [(5'h10):(1'h0)] reg553 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg552 = (1'h0);
  reg [(2'h2):(1'h0)] reg551 = (1'h0);
  reg [(5'h15):(1'h0)] reg550 = (1'h0);
  reg [(4'he):(1'h0)] reg549 = (1'h0);
  reg [(5'h14):(1'h0)] reg548 = (1'h0);
  reg [(5'h10):(1'h0)] reg547 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg546 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg545 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg544 = (1'h0);
  reg [(5'h15):(1'h0)] forvar543 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg542 = (1'h0);
  reg [(4'h8):(1'h0)] reg541 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg540 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg539 = (1'h0);
  reg [(4'ha):(1'h0)] reg538 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar537 = (1'h0);
  reg [(2'h3):(1'h0)] reg536 = (1'h0);
  reg [(3'h6):(1'h0)] reg535 = (1'h0);
  reg [(2'h3):(1'h0)] reg534 = (1'h0);
  reg [(5'h12):(1'h0)] reg533 = (1'h0);
  reg [(4'ha):(1'h0)] forvar532 = (1'h0);
  reg [(4'ha):(1'h0)] reg531 = (1'h0);
  reg [(5'h14):(1'h0)] forvar530 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg529 = (1'h0);
  reg [(4'he):(1'h0)] reg528 = (1'h0);
  reg [(4'h8):(1'h0)] reg527 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar526 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg525 = (1'h0);
  reg [(3'h6):(1'h0)] reg524 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg523 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg522 = (1'h0);
  reg [(5'h10):(1'h0)] reg521 = (1'h0);
  reg [(3'h4):(1'h0)] reg520 = (1'h0);
  reg [(3'h7):(1'h0)] forvar519 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg518 = (1'h0);
  reg [(3'h4):(1'h0)] reg517 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar516 = (1'h0);
  assign y = {wire639,
                 wire638,
                 wire637,
                 wire636,
                 wire635,
                 wire634,
                 wire633,
                 wire632,
                 wire631,
                 reg630,
                 reg629,
                 reg628,
                 forvar627,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 reg621,
                 reg620,
                 forvar619,
                 forvar618,
                 reg614,
                 reg617,
                 reg616,
                 reg615,
                 forvar614,
                 reg613,
                 reg612,
                 forvar611,
                 reg610,
                 forvar609,
                 reg608,
                 reg607,
                 wire606,
                 wire605,
                 reg604,
                 reg603,
                 reg602,
                 reg601,
                 reg600,
                 forvar595,
                 forvar591,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 reg588,
                 reg587,
                 forvar586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 reg580,
                 forvar579,
                 wire578,
                 wire577,
                 forvar569,
                 reg576,
                 reg575,
                 reg574,
                 reg573,
                 forvar572,
                 reg571,
                 reg570,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 forvar565,
                 reg564,
                 reg563,
                 reg562,
                 forvar561,
                 reg560,
                 reg559,
                 reg558,
                 wire557,
                 reg556,
                 reg555,
                 reg554,
                 reg553,
                 reg552,
                 reg551,
                 reg550,
                 reg549,
                 reg548,
                 reg547,
                 reg546,
                 reg545,
                 reg544,
                 forvar543,
                 reg542,
                 reg541,
                 reg540,
                 reg539,
                 reg538,
                 forvar537,
                 reg536,
                 reg535,
                 reg534,
                 reg533,
                 forvar532,
                 reg531,
                 forvar530,
                 reg529,
                 reg528,
                 reg527,
                 forvar526,
                 reg525,
                 reg524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 forvar519,
                 reg518,
                 reg517,
                 forvar516,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar516 = (1'h0); (forvar516 < (3'h4)); forvar516 = (forvar516 + (1'h1)))
        begin
          reg517 = ((({wire513,
                  (wire513 <<< wire515)} > wire515[(1'h1):(1'h0)]) ^ (^~(~^$unsigned(forvar516)))) ?
              $signed(forvar516[(1'h0):(1'h0)]) : ((((~(8'ha9)) ?
                      {wire513} : $unsigned((8'hb8))) ?
                  (wire515 ?
                      (forvar516 | wire514) : (wire512 < wire511)) : wire515[(2'h3):(1'h1)]) <<< {$signed(wire513[(3'h6):(1'h0)])}));
          reg518 <= $signed(wire515);
          for (forvar519 = (1'h0); (forvar519 < (1'h0)); forvar519 = (forvar519 + (1'h1)))
            begin
              reg520 <= $unsigned({($signed($unsigned(reg517)) ?
                      wire513 : ((-wire515) - (8'hbe)))});
              reg521 <= (~^$unsigned((forvar519[(3'h6):(3'h4)] ?
                  ($signed(wire513) != $signed(reg517)) : wire511)));
              reg522 <= ($unsigned((forvar516 ?
                  $unsigned((forvar519 ^ reg518)) : wire511)) ~^ (&$signed(wire513[(1'h0):(1'h0)])));
              reg523 <= wire514;
            end
        end
    end
  always
    @(posedge clk) begin
      reg524 <= {$signed(wire512)};
      reg525 <= $unsigned({(wire512 ?
              wire512[(1'h1):(1'h1)] : $signed(((8'ha6) ?
                  forvar519 : wire515))),
          $signed($signed((wire511 >> wire511)))});
    end
  always
    @(posedge clk) begin
      for (forvar526 = (1'h0); (forvar526 < (3'h4)); forvar526 = (forvar526 + (1'h1)))
        begin
          reg527 <= reg518[(2'h2):(2'h2)];
          reg528 <= (-$signed({$signed((~(8'haa)))}));
        end
      reg529 = $signed($unsigned(wire513));
      for (forvar530 = (1'h0); (forvar530 < (1'h1)); forvar530 = (forvar530 + (1'h1)))
        begin
          reg531 <= ((~&reg523[(2'h2):(2'h2)]) ^~ "xfwlFA8YIAGushcKeX5v");
          for (forvar532 = (1'h0); (forvar532 < (2'h2)); forvar532 = (forvar532 + (1'h1)))
            begin
              reg533 <= $unsigned((forvar516[(1'h0):(1'h0)] && $unsigned((^~reg522[(1'h1):(1'h0)]))));
              reg534 = (reg518 ?
                  ((reg525[(4'hb):(3'h7)] ?
                      $unsigned($signed(wire514)) : (forvar516[(1'h0):(1'h0)] || forvar530)) > forvar532[(2'h3):(2'h3)]) : $signed((reg529 + forvar519)));
              reg535 = $signed("CfutF1zUbuHr2Hmr37");
              reg536 <= $unsigned((($signed($signed(wire513)) <<< (reg531 ?
                  $signed((8'ha4)) : (~|reg520))) | (|(((8'hb1) | (8'hb6)) ?
                  reg531[(1'h0):(1'h0)] : reg534))));
            end
          for (forvar537 = (1'h0); (forvar537 < (3'h4)); forvar537 = (forvar537 + (1'h1)))
            begin
              reg538 = (reg535 ?
                  forvar516[(1'h0):(1'h0)] : (&((~$signed(reg527)) > forvar516)));
              reg539 = ($unsigned(reg520) == {$signed((&(reg528 ?
                      reg522 : forvar519)))});
              reg540 <= ({($signed((wire511 <<< reg522)) ?
                      (wire514[(3'h5):(1'h0)] + $unsigned(forvar519)) : $unsigned(reg523[(3'h4):(2'h2)])),
                  ("iqRDAG4ll" ?
                      (^~(reg535 >>> reg528)) : "EFDKk48Qe")} >>> $signed(reg522));
            end
          reg541 = (8'hab);
          reg542 = $unsigned(($unsigned($signed($signed(forvar526))) ?
              (~&{((8'hb5) ? reg524 : reg521),
                  wire511}) : $signed((wire515[(2'h3):(1'h1)] ?
                  $signed(reg517) : (wire511 >= (8'h9c))))));
        end
      if (reg539)
        begin
          for (forvar543 = (1'h0); (forvar543 < (1'h0)); forvar543 = (forvar543 + (1'h1)))
            begin
              reg544 = (~|forvar516[(1'h1):(1'h0)]);
              reg545 <= reg521[(3'h4):(2'h2)];
              reg546 <= ($signed($signed($unsigned($signed(reg539)))) ?
                  $unsigned(forvar532[(3'h5):(3'h4)]) : $signed({((reg533 ?
                              (8'hae) : reg524) ?
                          {wire512, reg535} : $unsigned(reg544)),
                      ((reg533 ? reg525 : (8'h9c)) ?
                          (reg534 <<< (8'haf)) : $signed(wire512))}));
              reg547 = reg517[(2'h3):(1'h1)];
            end
          if (($signed(reg539[(3'h4):(2'h2)]) ?
              (reg534[(1'h1):(1'h0)] + $unsigned(((~|reg520) ?
                  ((8'hb9) ?
                      wire513 : reg527) : $unsigned(reg525)))) : (-reg544[(2'h2):(1'h1)])))
            begin
              reg548 <= (reg540 != (8'haf));
              reg549 <= {"mDWGTEXKEMC"};
              reg550 = $signed({$unsigned(($unsigned(reg520) ?
                      $unsigned(reg523) : {reg533})),
                  ((~|(reg528 >= reg527)) ? $signed(reg541) : reg536)});
              reg551 <= (reg517 >= reg531[(3'h5):(2'h2)]);
            end
          else
            begin
              reg548 <= $signed(((reg540 ?
                      ($signed(reg527) ^~ (reg522 | forvar526)) : (reg538[(3'h4):(2'h2)] ?
                          {(8'hb8)} : reg538)) ?
                  (^~(!(reg518 != forvar537))) : ((forvar526 - (reg538 + wire515)) + $unsigned($signed(reg538)))));
              reg549 <= $signed(wire515);
              reg550 <= ("hmsF" <<< (~(((~|forvar530) >>> reg542[(2'h2):(1'h1)]) ?
                  ((reg544 >> reg535) < (reg534 ?
                      reg548 : reg549)) : ($signed(reg550) ?
                      (+(8'ha4)) : (8'ha0)))));
            end
          if ($signed($signed((8'hb4))))
            begin
              reg552 <= (((~&$signed((reg524 ? forvar516 : (8'ha5)))) ?
                      $signed({$unsigned((8'hb7)),
                          (reg529 ?
                              reg527 : reg536)}) : reg538[(2'h3):(1'h0)]) ?
                  (~$unsigned($unsigned($unsigned(wire514)))) : reg540);
              reg553 = forvar526[(1'h0):(1'h0)];
              reg554 = {reg538[(4'h8):(2'h2)],
                  $unsigned($signed($unsigned($unsigned(reg545))))};
              reg555 = wire514;
            end
          else
            begin
              reg552 = ({(reg535 - reg550)} && $signed("5ybha9laU"));
              reg553 <= (reg547 ~^ (8'ha3));
              reg554 <= ($signed(forvar537[(1'h1):(1'h0)]) - reg520[(2'h2):(1'h0)]);
            end
        end
      else
        begin
          for (forvar543 = (1'h0); (forvar543 < (3'h4)); forvar543 = (forvar543 + (1'h1)))
            begin
              reg544 = (^~((8'ha0) ~^ (~(~|reg517))));
              reg545 <= $signed(reg547[(4'h9):(3'h7)]);
              reg546 <= reg540;
              reg547 <= ($signed(($signed("1Sq") > reg555[(3'h4):(2'h3)])) ^ $signed($unsigned(reg549[(4'ha):(4'ha)])));
              reg548 <= $unsigned(($signed(reg521) ?
                  ($signed((~&reg542)) ?
                      (^(reg538 ?
                          forvar519 : (8'hbc))) : "kvNXoOgwMZPe") : reg534[(2'h3):(2'h3)]));
            end
        end
      reg556 <= $unsigned($signed($signed(reg527[(3'h7):(3'h5)])));
    end
  assign wire557 = reg542[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      reg558 <= forvar526[(3'h5):(3'h4)];
      if ("2RHFc5BX6Umx6XOx")
        begin
          reg559 <= forvar537;
          reg560 <= $signed(reg534[(2'h3):(1'h1)]);
          for (forvar561 = (1'h0); (forvar561 < (2'h3)); forvar561 = (forvar561 + (1'h1)))
            begin
              reg562 = $unsigned((~&$unsigned(($unsigned((8'ha5)) * (reg547 ?
                  reg518 : reg559)))));
              reg563 <= $signed({(&($signed(forvar537) >= reg559[(4'h9):(3'h4)]))});
            end
          reg564 <= ({(-(!reg559)),
              {$unsigned(reg551)}} || forvar532[(1'h1):(1'h0)]);
          for (forvar565 = (1'h0); (forvar565 < (2'h3)); forvar565 = (forvar565 + (1'h1)))
            begin
              reg566 <= reg562[(1'h1):(1'h1)];
              reg567 = (!$unsigned($unsigned({reg545[(3'h4):(1'h0)], reg550})));
              reg568 <= ((8'h9d) ?
                  ($unsigned(reg566) ?
                      (((reg544 ~^ reg542) ?
                          {(8'hb9)} : $unsigned((8'h9f))) > ($unsigned((8'ha9)) >>> wire557[(5'h10):(3'h6)])) : $signed($signed($signed(reg558)))) : $signed(((reg549 ?
                          $unsigned(forvar526) : $unsigned(reg535)) ?
                      $signed((reg564 ? reg559 : reg528)) : ($unsigned(reg560) ?
                          $signed(reg567) : (reg540 >>> reg552)))));
            end
        end
      else
        begin
          reg559 <= ($signed(reg531[(4'ha):(2'h3)]) ?
              (($signed($unsigned(reg554)) == $signed(wire557[(5'h13):(3'h4)])) > $unsigned($unsigned("hv"))) : ((~&($signed(forvar516) ?
                      "MkhpU0J" : $unsigned((8'h9e)))) ?
                  reg562[(2'h2):(1'h1)] : (+reg540)));
          reg560 = ($unsigned(((~&$unsigned(reg524)) >>> $unsigned((forvar526 ~^ reg535)))) ?
              "zDozE48hOSnH" : ("R89qouyUU049rRLIQlP" <= ($unsigned((~^(8'hbd))) >> ($signed(reg541) ?
                  $unsigned(reg542) : wire515))));
          for (forvar561 = (1'h0); (forvar561 < (2'h3)); forvar561 = (forvar561 + (1'h1)))
            begin
              reg562 = reg522;
            end
        end
      if (reg546[(3'h6):(3'h5)])
        begin
          reg569 = {{{((~wire513) ? (wire512 ? reg520 : reg518) : (8'hbe))}},
              reg523};
          reg570 = (reg533[(5'h12):(4'ha)] || (8'hb3));
          reg571 <= $signed(reg534[(2'h3):(2'h3)]);
          for (forvar572 = (1'h0); (forvar572 < (2'h3)); forvar572 = (forvar572 + (1'h1)))
            begin
              reg573 <= "LS";
              reg574 = $unsigned((reg541[(2'h3):(2'h2)] ?
                  $signed((~(|reg545))) : reg569[(3'h5):(1'h0)]));
              reg575 = reg548;
              reg576 <= (($signed(((-wire512) ? forvar537 : {reg518})) ?
                      ($unsigned($signed(reg541)) ?
                          $signed(forvar530[(5'h12):(5'h12)]) : {(reg544 ?
                                  (8'ha1) : reg545)}) : ((((8'h9f) ?
                                  forvar537 : reg566) ?
                              reg553[(4'hf):(3'h7)] : (8'hb0)) ?
                          $signed(reg574[(1'h0):(1'h0)]) : (forvar565[(5'h15):(2'h2)] != reg536[(2'h2):(2'h2)]))) ?
                  {(($unsigned(forvar516) >= $unsigned(reg539)) >> ($unsigned(reg563) ?
                          $signed(reg571) : forvar565[(5'h10):(4'hd)]))} : $signed(reg551[(2'h2):(1'h0)]));
            end
        end
      else
        begin
          for (forvar569 = (1'h0); (forvar569 < (2'h3)); forvar569 = (forvar569 + (1'h1)))
            begin
              reg570 = {($unsigned($unsigned((reg541 + forvar516))) >>> $unsigned(((reg539 ?
                      reg558 : (8'hba)) >>> (reg560 >> reg575))))};
              reg571 <= (reg569 >>> $unsigned(forvar537[(3'h4):(2'h2)]));
            end
        end
    end
  assign wire577 = wire514;
  assign wire578 = ((wire514[(1'h0):(1'h0)] ~^ {(8'had)}) ?
                       reg558[(4'h8):(3'h5)] : $unsigned((reg570[(1'h0):(1'h0)] ?
                           (~&forvar565[(2'h2):(1'h0)]) : ($unsigned(reg563) ?
                               forvar543 : reg551))));
  always
    @(posedge clk) begin
      for (forvar579 = (1'h0); (forvar579 < (1'h0)); forvar579 = (forvar579 + (1'h1)))
        begin
          if ($signed($unsigned({{$signed(reg550)}})))
            begin
              reg580 <= $unsigned((forvar561[(1'h1):(1'h1)] ?
                  $unsigned(reg540[(3'h4):(1'h0)]) : $unsigned($signed((reg566 ?
                      reg564 : reg563)))));
              reg581 <= reg569;
              reg582 <= $signed((~(!reg520)));
              reg583 <= (8'hb6);
              reg584 <= (8'hb3);
            end
          else
            begin
              reg580 <= (-(reg559 && (reg548 && (reg567[(1'h1):(1'h0)] ^ (forvar572 ?
                  reg554 : reg542)))));
              reg581 = $unsigned((8'ha1));
              reg582 <= $unsigned($unsigned((~|$unsigned(reg567[(2'h2):(1'h1)]))));
            end
          reg585 <= ((({reg571[(4'hc):(3'h4)]} ?
              "pVkyW0OPQFbXyewZ" : ($signed(reg548) ?
                  reg582[(4'hd):(4'hb)] : {(8'ha5)})) && forvar516) + $signed($unsigned((8'ha3))));
          for (forvar586 = (1'h0); (forvar586 < (2'h2)); forvar586 = (forvar586 + (1'h1)))
            begin
              reg587 = ($signed({forvar572}) ?
                  reg566 : (!(-reg551[(1'h0):(1'h0)])));
              reg588 <= ($unsigned(forvar565) > (((+{reg562}) > "VPsrox3pMZsEa3ErDQX7") ?
                  reg570[(4'hd):(2'h3)] : forvar561[(1'h0):(1'h0)]));
              reg589 <= reg546[(4'h9):(2'h3)];
            end
        end
      reg590 <= $signed((^~$unsigned(reg529)));
      if (($unsigned($unsigned(($signed(forvar586) ?
          $unsigned(wire512) : "ykERW3zU"))) == $unsigned($signed(reg580[(2'h3):(1'h1)]))))
        begin
          if ($signed(((8'ha5) != $unsigned($signed((-(7'h43)))))))
            begin
              reg591 = $unsigned(reg582[(4'hf):(4'h8)]);
              reg592 = reg556[(5'h12):(4'he)];
              reg593 <= reg566;
              reg594 <= {{reg574[(2'h2):(2'h2)]}};
            end
          else
            begin
              reg591 = $unsigned("bphQHBOsvqK9xx5N0");
              reg592 = reg552;
            end
          reg595 = forvar586;
          if (({reg542[(1'h1):(1'h0)],
              (~&reg563)} + ((((-reg541) && ((8'hbf) > reg594)) != (-(reg528 ?
              (8'hbc) : reg582))) < ($unsigned(((8'hbe) ^~ forvar565)) ?
              ($unsigned((7'h43)) ^~ forvar519[(1'h0):(1'h0)]) : (|(|reg522))))))
            begin
              reg596 = $unsigned($signed(reg568));
              reg597 = ((((~|reg560[(4'hd):(3'h4)]) ?
                      (forvar543[(5'h13):(4'he)] < reg573[(3'h7):(1'h1)]) : ((reg575 >>> reg576) + reg595[(2'h3):(2'h3)])) ?
                  $signed((~&(reg539 ? wire577 : forvar530))) : (-(+((8'hbf) ?
                      (8'ha1) : reg567)))) && ($signed(((reg555 ?
                  reg535 : reg527) <<< reg570)) << $signed((~^(~|reg563)))));
            end
          else
            begin
              reg596 <= $unsigned((reg596[(3'h6):(2'h3)] ?
                  $unsigned(($unsigned(wire514) ?
                      $signed(forvar526) : $unsigned(forvar516))) : {{(~^reg547),
                          $signed(reg553)},
                      $unsigned($unsigned(reg523))}));
              reg597 <= $signed(reg570);
              reg598 <= (^~$unsigned({$signed((reg580 ? reg574 : reg570)),
                  reg589[(2'h2):(1'h1)]}));
              reg599 <= ($unsigned(forvar519[(2'h3):(2'h2)]) ^~ reg585);
            end
        end
      else
        begin
          for (forvar591 = (1'h0); (forvar591 < (2'h2)); forvar591 = (forvar591 + (1'h1)))
            begin
              reg592 <= "MQT";
              reg593 <= (8'hb3);
              reg594 <= {{(reg555[(3'h7):(3'h7)] ?
                          $signed((reg528 && reg566)) : forvar537[(3'h4):(1'h1)])}};
            end
          for (forvar595 = (1'h0); (forvar595 < (2'h3)); forvar595 = (forvar595 + (1'h1)))
            begin
              reg596 = {$signed($signed($unsigned($signed(reg564))))};
              reg597 <= ((({(^~forvar516), wire512} ?
                  $signed({reg574}) : (reg583[(5'h10):(1'h0)] - {reg538})) <<< $signed(reg536)) | reg540[(4'hc):(4'h8)]);
              reg598 <= $signed(reg576);
            end
          if ((~|(~|$unsigned({(+wire515), $unsigned(reg574)}))))
            begin
              reg599 = reg588[(4'hd):(4'ha)];
              reg600 <= ((8'hb9) ?
                  (("oZQHRTMOXw9eCPtm" && {(reg521 ?
                          reg595 : reg518)}) >= reg567) : (^~reg593));
              reg601 = reg536[(2'h2):(1'h1)];
              reg602 <= reg584[(4'ha):(4'h8)];
            end
          else
            begin
              reg599 = ($signed(reg554) > ((^~$signed(reg544)) + {$unsigned($unsigned(reg575))}));
              reg600 = ({$unsigned({$signed(reg570)}),
                      (|(&reg539[(3'h5):(3'h4)]))} ?
                  $unsigned(forvar530[(4'hf):(4'hf)]) : {reg520, forvar537});
              reg601 = $signed(reg588);
              reg602 = $signed(reg553[(4'he):(4'he)]);
              reg603 = {(((reg567[(1'h0):(1'h0)] ?
                      reg541[(3'h6):(3'h4)] : $unsigned(reg520)) | $unsigned(reg549)) >= (+(!$unsigned(wire513)))),
                  $unsigned(forvar561)};
            end
        end
      reg604 = ((reg548 + wire577[(1'h0):(1'h0)]) ?
          forvar591 : forvar565[(5'h13):(1'h1)]);
    end
  assign wire605 = (~^$unsigned((8'h9c)));
  assign wire606 = $signed(reg587);
  always
    @(posedge clk) begin
      reg607 = "nF";
      reg608 = (reg581[(3'h5):(3'h4)] ~^ $signed(wire514[(2'h3):(1'h1)]));
      for (forvar609 = (1'h0); (forvar609 < (1'h1)); forvar609 = (forvar609 + (1'h1)))
        begin
          reg610 <= reg574;
          for (forvar611 = (1'h0); (forvar611 < (3'h4)); forvar611 = (forvar611 + (1'h1)))
            begin
              reg612 <= $unsigned($unsigned(($unsigned({(8'ha8)}) ?
                  $signed($signed(reg554)) : ((wire606 ? reg607 : reg520) ?
                      (~|reg576) : {reg545, reg587}))));
              reg613 = reg599;
            end
        end
      if ($signed($unsigned((7'h43))))
        begin
          for (forvar614 = (1'h0); (forvar614 < (2'h3)); forvar614 = (forvar614 + (1'h1)))
            begin
              reg615 <= reg539;
              reg616 = $signed($unsigned({wire511[(3'h6):(1'h1)]}));
              reg617 <= ({$unsigned(((8'hac) < reg541)),
                      $unsigned(({reg536, (8'hb6)} < reg535[(1'h0):(1'h0)]))} ?
                  forvar516 : (($unsigned((forvar611 | wire514)) ?
                          $unsigned((wire605 ?
                              reg580 : reg529)) : $unsigned((!(8'ha1)))) ?
                      (reg540 ?
                          forvar537 : forvar543[(4'hc):(4'hc)]) : (8'haa)));
            end
        end
      else
        begin
          reg614 <= forvar530[(2'h3):(1'h1)];
          reg615 <= reg581;
          reg616 <= $signed($signed($unsigned({(~|reg549),
              $unsigned(reg548)})));
        end
      for (forvar618 = (1'h0); (forvar618 < (1'h1)); forvar618 = (forvar618 + (1'h1)))
        begin
          for (forvar619 = (1'h0); (forvar619 < (2'h2)); forvar619 = (forvar619 + (1'h1)))
            begin
              reg620 = (~(^$unsigned($signed((forvar586 ? reg584 : reg522)))));
              reg621 <= $signed($unsigned({$signed(reg533), reg566}));
            end
          if (reg556)
            begin
              reg622 = ((8'h9d) >>> ({$unsigned((reg594 ? reg575 : reg523)),
                      ((8'hb4) * (-reg558))} ?
                  reg620 : (((8'hbf) <= {wire512}) > ((wire515 & reg539) > (reg590 ?
                      forvar579 : (7'h44))))));
              reg623 <= (-$signed(($signed($unsigned(reg582)) - wire512[(1'h1):(1'h0)])));
              reg624 <= ($unsigned((reg601[(1'h0):(1'h0)] ?
                      $unsigned((~|reg539)) : $unsigned($signed(forvar532)))) ?
                  $unsigned(reg531[(3'h6):(2'h2)]) : $unsigned(reg604[(2'h3):(1'h0)]));
              reg625 <= $unsigned($signed((~$signed((forvar519 > (8'hbb))))));
            end
          else
            begin
              reg622 <= reg517[(2'h2):(2'h2)];
              reg623 = (reg521[(4'hc):(1'h0)] ?
                  (~|$signed(forvar516[(2'h2):(1'h0)])) : (8'ha1));
              reg624 = (!($signed(((reg560 ? reg542 : (8'h9e)) ?
                  reg582[(2'h2):(1'h0)] : (|(8'hb9)))) - (forvar516[(1'h1):(1'h0)] ?
                  $unsigned(reg525[(4'ha):(3'h6)]) : $signed($unsigned(reg608)))));
              reg625 = ((($unsigned((!reg531)) == ($signed(forvar537) - {(8'hb4),
                      reg552})) ?
                  $unsigned((forvar569[(4'hf):(3'h4)] ?
                      reg616 : (8'ha3))) : (($signed((8'hb0)) & forvar532[(4'ha):(3'h6)]) < $unsigned({wire578}))) > ($signed(reg538[(3'h7):(3'h4)]) + (((reg553 ^ reg527) <= (reg523 ?
                      reg599 : forvar595)) ?
                  {(~reg584)} : (8'h9e))));
            end
          reg626 = $unsigned(forvar579);
          for (forvar627 = (1'h0); (forvar627 < (1'h1)); forvar627 = (forvar627 + (1'h1)))
            begin
              reg628 <= $signed(reg602[(3'h7):(2'h3)]);
              reg629 = (+reg602);
              reg630 <= reg540;
            end
        end
    end
  assign wire631 = $unsigned(((((~^reg539) ?
                               (reg520 >>> reg521) : (reg599 ?
                                   forvar565 : reg541)) ?
                           $unsigned((-(8'hbc))) : $signed(reg549[(4'h9):(3'h6)])) ?
                       forvar569[(2'h3):(1'h1)] : (^~{(forvar519 ?
                               reg602 : reg547)})));
  assign wire632 = $signed(reg574[(5'h14):(5'h14)]);
  assign wire633 = reg529;
  assign wire634 = forvar579;
  assign wire635 = (8'hac);
  assign wire636 = $unsigned($unsigned($signed(($signed((8'h9e)) ?
                       reg548[(4'hd):(3'h4)] : (reg608 || reg546)))));
  assign wire637 = (8'hb2);
  assign wire638 = (forvar569 ?
                       (wire636 ?
                           (~|(8'hac)) : (7'h41)) : (reg559[(4'ha):(3'h7)] ?
                           ($signed($unsigned(forvar586)) ?
                               ((^~reg599) & reg523) : (7'h40)) : $signed(reg548[(1'h0):(1'h0)])));
  assign wire639 = $unsigned(reg552[(3'h6):(3'h6)]);
endmodule