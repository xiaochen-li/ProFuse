(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire4, wire3, wire2, wire1, wire0);
  output wire [(32'h40f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire4;
  input wire [(4'hf):(1'h0)] wire3;
  input wire [(5'h12):(1'h0)] wire2;
  input wire [(5'h16):(1'h0)] wire1;
  input wire signed [(4'h9):(1'h0)] wire0;
  wire [(3'h5):(1'h0)] wire1771;
  wire signed [(5'h13):(1'h0)] wire1769;
  wire signed [(2'h2):(1'h0)] wire1768;
  wire [(5'h14):(1'h0)] wire1745;
  wire [(4'hb):(1'h0)] wire1744;
  wire [(4'ha):(1'h0)] wire1740;
  wire signed [(5'h12):(1'h0)] wire52;
  wire signed [(5'h15):(1'h0)] wire38;
  wire signed [(5'h16):(1'h0)] wire37;
  wire signed [(2'h2):(1'h0)] wire35;
  wire signed [(5'h17):(1'h0)] wire8;
  wire signed [(5'h11):(1'h0)] wire7;
  reg [(4'hb):(1'h0)] reg1767 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1765 = (1'h0);
  reg [(3'h7):(1'h0)] reg1761 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1755 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1754 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1751 = (1'h0);
  reg [(4'h9):(1'h0)] reg1749 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1746 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1743 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg10 = (1'h0);
  reg [(3'h6):(1'h0)] reg13 = (1'h0);
  reg [(4'hd):(1'h0)] reg14 = (1'h0);
  reg [(4'h9):(1'h0)] reg15 = (1'h0);
  reg [(5'h10):(1'h0)] reg17 = (1'h0);
  reg [(2'h2):(1'h0)] reg18 = (1'h0);
  reg [(4'ha):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg23 = (1'h0);
  reg [(4'ha):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg25 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg26 = (1'h0);
  reg [(5'h13):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg29 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg36 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg39 = (1'h0);
  reg [(5'h11):(1'h0)] reg41 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg47 = (1'h0);
  reg [(5'h17):(1'h0)] reg49 = (1'h0);
  reg [(5'h14):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg51 = (1'h0);
  reg [(5'h10):(1'h0)] reg1766 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1764 = (1'h0);
  reg [(3'h7):(1'h0)] reg1763 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1762 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1760 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1759 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1758 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1747 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1757 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1756 = (1'h0);
  reg [(5'h11):(1'h0)] reg1753 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1752 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1750 = (1'h0);
  reg [(5'h13):(1'h0)] reg1748 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1747 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1742 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg48 = (1'h0);
  reg [(3'h5):(1'h0)] reg46 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg45 = (1'h0);
  reg [(3'h7):(1'h0)] reg44 = (1'h0);
  reg [(4'h8):(1'h0)] reg43 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg42 = (1'h0);
  reg [(4'hc):(1'h0)] reg40 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg34 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg33 = (1'h0);
  reg [(2'h3):(1'h0)] reg32 = (1'h0);
  reg [(3'h7):(1'h0)] reg31 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg28 = (1'h0);
  reg [(2'h3):(1'h0)] reg22 = (1'h0);
  reg [(5'h10):(1'h0)] reg20 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg19 = (1'h0);
  reg [(2'h3):(1'h0)] reg16 = (1'h0);
  reg [(4'ha):(1'h0)] forvar12 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg11 = (1'h0);
  reg [(3'h4):(1'h0)] forvar9 = (1'h0);
  reg [(3'h4):(1'h0)] reg6 = (1'h0);
  reg [(3'h7):(1'h0)] forvar5 = (1'h0);
  assign y = {wire1771,
                 wire1769,
                 wire1768,
                 wire1745,
                 wire1744,
                 wire1740,
                 wire52,
                 wire38,
                 wire37,
                 wire35,
                 wire8,
                 wire7,
                 reg1767,
                 reg1765,
                 reg1761,
                 reg1755,
                 reg1754,
                 reg1751,
                 reg1749,
                 reg1746,
                 reg1743,
                 reg10,
                 reg13,
                 reg14,
                 reg15,
                 reg17,
                 reg18,
                 reg21,
                 reg23,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 reg29,
                 reg30,
                 reg36,
                 reg39,
                 reg41,
                 reg47,
                 reg49,
                 reg50,
                 reg51,
                 reg1766,
                 forvar1764,
                 reg1763,
                 reg1762,
                 reg1760,
                 reg1759,
                 forvar1758,
                 reg1747,
                 reg1757,
                 reg1756,
                 reg1753,
                 reg1752,
                 reg1750,
                 reg1748,
                 forvar1747,
                 reg1742,
                 reg48,
                 reg46,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg40,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg28,
                 reg22,
                 reg20,
                 reg19,
                 reg16,
                 forvar12,
                 reg11,
                 forvar9,
                 reg6,
                 forvar5,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar5 = (1'h0); (forvar5 < (3'h4)); forvar5 = (forvar5 + (1'h1)))
        begin
          reg6 = $unsigned(((~&(~|(wire0 ?
              wire1 : wire0))) <= wire4[(4'hc):(4'hb)]));
        end
    end
  assign wire7 = {((({wire3} - $signed(wire0)) << ((8'hae) ?
                         wire1[(4'ha):(4'h9)] : wire4[(2'h3):(2'h3)])) ~^ (^((wire4 + wire3) > (8'hb4))))};
  assign wire8 = {wire7,
                     (^(($unsigned(wire4) ?
                             (wire1 >= wire7) : ((7'h41) ^~ wire2)) ?
                         (wire1 - ((7'h44) ?
                             wire2 : wire4)) : ($unsigned(wire4) ?
                             ((8'hb6) ? wire0 : wire2) : (wire3 ?
                                 wire1 : wire4))))};
  always
    @(posedge clk) begin
      for (forvar9 = (1'h0); (forvar9 < (3'h4)); forvar9 = (forvar9 + (1'h1)))
        begin
          reg10 <= $signed((!(wire4 ? $signed($unsigned(wire4)) : (8'ha3))));
          reg11 = wire4;
        end
      if (wire3[(3'h6):(1'h0)])
        begin
          for (forvar12 = (1'h0); (forvar12 < (1'h1)); forvar12 = (forvar12 + (1'h1)))
            begin
              reg13 <= (7'h43);
              reg14 <= wire0;
              reg15 <= wire7;
            end
          reg16 = (|$signed(forvar12[(3'h7):(3'h5)]));
          reg17 <= $signed((^~$unsigned(wire0)));
          reg18 <= $unsigned(wire1[(5'h16):(4'ha)]);
        end
      else
        begin
          for (forvar12 = (1'h0); (forvar12 < (2'h2)); forvar12 = (forvar12 + (1'h1)))
            begin
              reg13 <= $unsigned($unsigned($unsigned($signed((wire1 ?
                  forvar9 : (8'hab))))));
            end
        end
      if (wire1[(4'h9):(4'h8)])
        begin
          reg19 = reg15[(1'h0):(1'h0)];
          reg20 = (~^reg17);
          if ($unsigned($unsigned(((reg13 > $signed((8'ha8))) ?
              ((reg13 ? reg20 : forvar12) >= reg13[(2'h3):(1'h1)]) : (reg11 ?
                  $signed(wire3) : (reg10 ? wire8 : reg17))))))
            begin
              reg21 <= reg19;
              reg22 = forvar9;
              reg23 <= $signed((~|(8'ha1)));
            end
          else
            begin
              reg21 <= reg13;
              reg23 <= (|(wire8[(1'h1):(1'h0)] ?
                  {$signed($signed(wire2)),
                      reg18[(1'h1):(1'h1)]} : $unsigned(reg13)));
              reg24 <= $signed((~&{wire7}));
              reg25 <= reg16;
              reg26 <= (-$signed($signed((!$signed((7'h48))))));
            end
          if (reg22[(2'h2):(2'h2)])
            begin
              reg27 <= ($unsigned(({(reg18 ? reg17 : (8'hb3))} <<< (~((8'h9f) ?
                      reg10 : reg22)))) ?
                  reg24 : $unsigned($unsigned((((8'h9c) ?
                      wire0 : wire7) - $unsigned(reg13)))));
              reg28 = (^~($signed({forvar12[(2'h2):(2'h2)]}) | forvar9));
              reg29 <= (wire2[(3'h7):(3'h7)] ?
                  (($unsigned(wire1) * $unsigned((wire3 ? reg10 : reg20))) ?
                      $signed(reg23) : (-wire8)) : (8'hb5));
            end
          else
            begin
              reg27 <= (~&($unsigned(wire3[(2'h2):(2'h2)]) <<< $unsigned($unsigned($signed(wire7)))));
              reg29 <= (^((reg13 > {reg17}) ?
                  reg26[(2'h3):(1'h0)] : (~|(~&(wire3 ? (8'ha2) : reg25)))));
              reg30 <= {reg26};
              reg31 = reg20[(3'h6):(1'h0)];
              reg32 = $unsigned((~($signed((~&(8'hb8))) << $signed((~^reg27)))));
            end
        end
      else
        begin
          if ({((reg24 <<< $unsigned((wire4 ? reg25 : reg31))) ?
                  reg14[(2'h3):(2'h2)] : $unsigned((reg18 * (reg21 || reg21)))),
              $signed($signed({reg27[(1'h0):(1'h0)],
                  (reg30 ? wire0 : reg10)}))})
            begin
              reg21 <= (($signed($unsigned((reg15 + forvar12))) >>> ((wire8[(2'h3):(1'h1)] == reg11[(1'h0):(1'h0)]) ?
                      ($unsigned(forvar9) ?
                          (reg16 ~^ (8'hb0)) : (^~reg18)) : reg19)) ?
                  ((((reg25 ? reg26 : reg25) ? $unsigned(reg15) : {wire0}) ?
                      $signed(reg26[(3'h6):(1'h0)]) : $unsigned((reg28 || reg25))) << (-wire1)) : (-reg19[(4'hb):(1'h1)]));
              reg22 = (^forvar12);
              reg23 <= wire8;
              reg24 <= (forvar12[(3'h5):(1'h1)] > (((8'hb0) << reg15[(3'h5):(3'h4)]) ^~ (-$signed($signed((8'hae))))));
              reg28 = (^~(($unsigned(reg27) || wire0[(3'h5):(1'h0)]) == $signed(reg29)));
            end
          else
            begin
              reg19 = (reg21 ?
                  $unsigned(($unsigned((wire4 + reg14)) > ($signed(reg18) ?
                      (reg14 ?
                          reg26 : reg17) : $signed(reg28)))) : reg17[(1'h0):(1'h0)]);
              reg20 = ((wire2[(4'hd):(4'h9)] < $unsigned(($unsigned(wire3) <= {reg22,
                      reg31}))) ?
                  (wire8 | $signed(reg10)) : ((((~forvar9) ?
                          (7'h40) : reg21[(3'h5):(2'h3)]) ?
                      reg28 : ($signed(reg28) ?
                          (^~forvar12) : (reg18 == (8'ha2)))) ^~ (~reg29)));
              reg22 = $signed((~&(reg26[(3'h5):(2'h2)] ?
                  reg20 : {(reg24 != reg20)})));
              reg23 <= $signed($unsigned($unsigned({$signed(reg17)})));
              reg28 = (&((+(~|reg23[(2'h3):(2'h3)])) ?
                  (((wire3 * reg15) * (wire3 ? reg31 : reg13)) ?
                      (8'hb6) : reg28) : wire4));
            end
        end
      reg33 = $signed(reg24);
    end
  always
    @(posedge clk) begin
      reg34 = $signed(($unsigned($signed({reg29, reg10})) ?
          reg18[(2'h2):(1'h1)] : $signed(wire4)));
    end
  assign wire35 = (!(^((7'h4a) >= ($unsigned(reg29) ~^ $signed(reg18)))));
  always
    @(posedge clk) begin
      reg36 <= (reg30 != $signed($signed((7'h42))));
    end
  assign wire37 = reg27;
  assign wire38 = $signed($unsigned(reg23[(2'h2):(1'h0)]));
  always
    @(posedge clk) begin
      reg39 <= $signed((!{((wire8 ? (8'hac) : reg15) ? reg36 : wire35),
          $unsigned({wire7, (8'hb7)})}));
      if ((7'h48))
        begin
          if (($signed(wire37) & wire1))
            begin
              reg40 = wire7[(4'ha):(1'h1)];
            end
          else
            begin
              reg41 <= reg14;
              reg42 = ((~$signed(reg17[(4'hb):(2'h3)])) | reg18);
              reg43 = ((-reg39[(2'h3):(2'h3)]) ?
                  reg13 : ((^~reg41[(4'hd):(1'h0)]) ?
                      ({(!reg39)} ?
                          ((7'h41) ?
                              $unsigned(reg27) : (wire7 ?
                                  wire8 : reg23)) : (reg27[(4'h9):(3'h5)] ?
                              (wire37 ? reg40 : wire0) : reg36)) : {(wire1 ?
                              (wire37 ? reg13 : reg30) : (~^reg26))}));
              reg44 = ($signed(reg29) ?
                  (7'h48) : (^~$unsigned((~^$signed((8'hb0))))));
              reg45 = $signed(reg27);
            end
          if (reg39)
            begin
              reg46 = reg42;
              reg47 <= wire3;
              reg48 = (reg21[(4'h8):(1'h1)] ?
                  ((({wire38} ?
                      {wire0} : {reg47}) <= reg40) >>> wire8) : $unsigned($signed((&(~(7'h48))))));
            end
          else
            begin
              reg47 <= (~&reg41);
              reg48 = reg15;
              reg49 <= (8'hb6);
              reg50 <= (reg47[(4'h8):(1'h1)] ?
                  reg44[(2'h2):(1'h0)] : reg41[(5'h11):(3'h7)]);
            end
        end
      else
        begin
          reg40 = $signed(wire7);
        end
    end
  always
    @(posedge clk) begin
      reg51 <= reg14[(4'hb):(4'h9)];
    end
  assign wire52 = (~&reg25);
  module53 #() modinst1741 (.y(wire1740), .wire57(reg24), .wire55(wire38), .wire54(reg17), .wire58(reg23), .wire56(wire2), .clk(clk));
  always
    @(posedge clk) begin
      reg1742 = $signed(reg49);
      reg1743 <= ($unsigned($signed(((^reg24) ?
          $unsigned(wire3) : {reg39}))) | reg30);
    end
  assign wire1744 = $unsigned($unsigned(((|(reg41 - reg30)) <= {reg29})));
  assign wire1745 = {wire37[(5'h16):(4'hd)],
                        (&$unsigned($unsigned((~&reg15))))};
  always
    @(posedge clk) begin
      reg1746 <= ($signed($signed($unsigned((reg30 ?
          wire1744 : wire1)))) >>> (reg27 * wire38[(5'h14):(2'h2)]));
    end
  always
    @(posedge clk) begin
      if ($signed((8'hbc)))
        begin
          for (forvar1747 = (1'h0); (forvar1747 < (2'h3)); forvar1747 = (forvar1747 + (1'h1)))
            begin
              reg1748 = $unsigned(((reg36[(2'h2):(2'h2)] & (|((7'h43) ?
                      reg49 : reg41))) ?
                  wire0 : (wire3[(3'h6):(2'h2)] ?
                      wire52[(4'hc):(1'h0)] : (reg14 ^~ {reg25}))));
              reg1749 <= (~(reg51 + ((reg47 ? (&reg29) : (reg21 < wire52)) ?
                  $unsigned((wire7 << (8'ha7))) : (8'ha7))));
            end
          reg1750 = (~^$signed($signed($signed($signed(wire8)))));
          if (((($unsigned((~^reg50)) != wire37) ?
              (~&((wire1744 & reg50) <<< wire2)) : $signed(wire3)) >> (8'hae)))
            begin
              reg1751 <= ($signed(wire0[(2'h2):(1'h1)]) >= ($unsigned(reg23) ?
                  (~&((reg36 ? reg15 : reg14) ?
                      $signed(wire35) : (reg23 ~^ (8'hb8)))) : ($signed({reg1748}) ^ ($signed(reg30) && reg10[(3'h4):(1'h0)]))));
              reg1752 = ((~|$unsigned(($unsigned(reg30) ?
                      (reg24 ? forvar1747 : reg14) : wire52[(4'hc):(1'h0)]))) ?
                  ((!($signed((8'hb4)) >= (-(8'ha1)))) && reg1743[(1'h1):(1'h1)]) : $unsigned({((+reg1749) ?
                          $signed(wire1740) : (wire0 ?
                              (8'hb1) : forvar1747))}));
              reg1753 = $signed((&({(|(8'h9d))} ?
                  $unsigned((7'h47)) : (~&reg39))));
              reg1754 <= $unsigned(reg41);
            end
          else
            begin
              reg1752 = reg1751[(2'h2):(1'h1)];
              reg1753 = {$signed(((wire7 ?
                      $unsigned(wire7) : {(8'hbd)}) < $unsigned($unsigned(reg41)))),
                  reg39[(2'h3):(1'h1)]};
              reg1754 <= $signed(reg47);
              reg1755 <= (-reg18);
            end
          reg1756 = ($unsigned(wire0[(2'h3):(2'h3)]) * wire1740);
          reg1757 = reg1752;
        end
      else
        begin
          reg1747 = ($signed($unsigned(((+reg36) ?
              $unsigned(reg1755) : reg1751))) >= (+reg1753));
          reg1748 = $unsigned(($signed(((+reg13) && (8'h9f))) ?
              $signed($signed((reg1750 ?
                  reg1755 : (8'had)))) : (reg1754[(4'hf):(1'h0)] ?
                  ((+(8'hbc)) >>> (^~reg1751)) : ($unsigned((8'haf)) ~^ $signed((8'hbe))))));
          reg1749 <= $signed((^~(((reg1756 << reg10) ?
              {reg1754} : reg1752) == $unsigned($unsigned(reg23)))));
          reg1751 <= (~&$unsigned((wire1740[(3'h6):(2'h3)] >= (-(8'hb1)))));
          reg1752 = $signed(($unsigned(((reg1757 ? (8'hb0) : reg30) ?
                  {reg1748} : wire8[(3'h4):(3'h4)])) ?
              reg1754 : (&reg25)));
        end
      for (forvar1758 = (1'h0); (forvar1758 < (3'h4)); forvar1758 = (forvar1758 + (1'h1)))
        begin
          if (wire1744[(4'hb):(1'h0)])
            begin
              reg1759 = $signed((reg1753[(3'h5):(2'h2)] + ((wire7 ?
                  (~^reg21) : (reg47 ^ (7'h45))) < (~^(reg15 ?
                  reg1751 : reg1752)))));
              reg1760 = $signed(reg1751[(2'h3):(1'h0)]);
              reg1761 <= ((8'ha2) << $signed($unsigned(($unsigned(wire8) ?
                  wire2[(2'h2):(1'h0)] : (reg50 ? reg1756 : (7'h45))))));
              reg1762 = $unsigned((|(reg14 >> reg27[(5'h12):(1'h1)])));
              reg1763 = reg1754[(5'h11):(4'he)];
            end
          else
            begin
              reg1759 = (&(&$unsigned(reg26)));
              reg1760 = $signed($unsigned($unsigned(reg1743)));
              reg1761 <= (wire1740 > reg27);
            end
          for (forvar1764 = (1'h0); (forvar1764 < (2'h2)); forvar1764 = (forvar1764 + (1'h1)))
            begin
              reg1765 <= {($unsigned($signed(reg1756[(3'h4):(2'h2)])) * $signed($signed($unsigned(reg30)))),
                  $signed($unsigned((7'h42)))};
              reg1766 = reg1746;
              reg1767 <= wire2;
            end
        end
    end
  assign wire1768 = {{(+$unsigned(wire35)),
                            (-((reg41 < reg1751) || $unsigned(reg23)))},
                        wire2[(4'h9):(4'h9)]};
  module937 #() modinst1770 (.wire940(reg49), .wire941(wire1), .y(wire1769), .clk(clk), .wire938(wire8), .wire939(reg51));
  assign wire1771 = ((~^$signed(({reg36, (8'ha8)} > (reg1743 ?
                            wire1745 : reg41)))) ?
                        (!((wire1744[(3'h7):(3'h6)] ?
                                $signed(wire2) : (^~(8'ha2))) ?
                            {$unsigned(wire3),
                                (wire35 < reg41)} : $unsigned($unsigned(reg15)))) : ((^{(wire37 + wire7),
                            (reg25 <<< reg30)}) == $signed(reg18[(2'h2):(1'h0)])));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module53  (y, clk, wire58, wire57, wire56, wire55, wire54);
  output wire [(32'h844):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire58;
  input wire [(4'ha):(1'h0)] wire57;
  input wire signed [(4'ha):(1'h0)] wire56;
  input wire signed [(5'h15):(1'h0)] wire55;
  input wire signed [(5'h10):(1'h0)] wire54;
  wire signed [(5'h13):(1'h0)] wire1685;
  wire signed [(3'h4):(1'h0)] wire1601;
  wire signed [(3'h6):(1'h0)] wire1599;
  wire [(4'hd):(1'h0)] wire659;
  wire [(5'h15):(1'h0)] wire70;
  wire signed [(4'hf):(1'h0)] wire1723;
  wire signed [(3'h5):(1'h0)] wire1724;
  wire [(3'h6):(1'h0)] wire1735;
  reg signed [(3'h7):(1'h0)] reg1739 = (1'h0);
  reg [(4'hb):(1'h0)] reg1738 = (1'h0);
  reg [(2'h2):(1'h0)] reg1734 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1730 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1729 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1727 = (1'h0);
  reg [(3'h4):(1'h0)] reg1720 = (1'h0);
  reg [(5'h16):(1'h0)] reg1719 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1718 = (1'h0);
  reg [(2'h2):(1'h0)] reg1716 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1715 = (1'h0);
  reg [(2'h3):(1'h0)] reg1713 = (1'h0);
  reg [(2'h2):(1'h0)] reg1712 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1710 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1709 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1706 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1705 = (1'h0);
  reg [(3'h5):(1'h0)] reg1704 = (1'h0);
  reg [(5'h16):(1'h0)] reg1702 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1701 = (1'h0);
  reg [(4'hd):(1'h0)] reg1700 = (1'h0);
  reg [(5'h11):(1'h0)] reg1699 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1696 = (1'h0);
  reg [(4'hb):(1'h0)] reg1695 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1689 = (1'h0);
  reg [(4'h9):(1'h0)] reg678 = (1'h0);
  reg [(4'ha):(1'h0)] reg675 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg672 = (1'h0);
  reg [(5'h17):(1'h0)] reg670 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg668 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg666 = (1'h0);
  reg [(4'ha):(1'h0)] reg664 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg663 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg661 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg68 = (1'h0);
  reg [(5'h15):(1'h0)] reg64 = (1'h0);
  reg [(3'h6):(1'h0)] reg63 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg61 = (1'h0);
  reg [(5'h13):(1'h0)] reg59 = (1'h0);
  reg [(3'h5):(1'h0)] reg1603 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1605 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1606 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1607 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1608 = (1'h0);
  reg [(5'h15):(1'h0)] reg1609 = (1'h0);
  reg [(4'h8):(1'h0)] reg1620 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1621 = (1'h0);
  reg [(4'hf):(1'h0)] reg1625 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1627 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1631 = (1'h0);
  reg [(4'hb):(1'h0)] reg1633 = (1'h0);
  reg [(4'h9):(1'h0)] reg1635 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1638 = (1'h0);
  reg [(4'hd):(1'h0)] reg1639 = (1'h0);
  reg [(3'h4):(1'h0)] reg1640 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1645 = (1'h0);
  reg [(3'h6):(1'h0)] reg1647 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1654 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1656 = (1'h0);
  reg [(4'hc):(1'h0)] reg1657 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1658 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1659 = (1'h0);
  reg [(5'h10):(1'h0)] reg1664 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1665 = (1'h0);
  reg [(4'hb):(1'h0)] reg1666 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1670 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1672 = (1'h0);
  reg [(5'h18):(1'h0)] reg1674 = (1'h0);
  reg [(4'hc):(1'h0)] reg1676 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1684 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1737 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1733 = (1'h0);
  reg [(4'he):(1'h0)] forvar1732 = (1'h0);
  reg [(4'h8):(1'h0)] reg1731 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1728 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1726 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1725 = (1'h0);
  reg [(5'h16):(1'h0)] reg1722 = (1'h0);
  reg [(5'h10):(1'h0)] reg1721 = (1'h0);
  reg [(5'h11):(1'h0)] reg1717 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1714 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1711 = (1'h0);
  reg [(3'h6):(1'h0)] reg1708 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1707 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1703 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1698 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1697 = (1'h0);
  reg [(5'h12):(1'h0)] reg1690 = (1'h0);
  reg [(3'h4):(1'h0)] reg1697 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1696 = (1'h0);
  reg [(4'hf):(1'h0)] reg1694 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1693 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1692 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1691 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1690 = (1'h0);
  reg [(5'h15):(1'h0)] reg1688 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1687 = (1'h0);
  reg [(5'h16):(1'h0)] reg1683 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1682 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1681 = (1'h0);
  reg [(3'h4):(1'h0)] reg1680 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1679 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1678 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1677 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1675 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1673 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1671 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1669 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1668 = (1'h0);
  reg [(5'h15):(1'h0)] reg1667 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1663 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1662 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1661 = (1'h0);
  reg [(5'h15):(1'h0)] reg1660 = (1'h0);
  reg [(5'h12):(1'h0)] reg1655 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1653 = (1'h0);
  reg [(5'h16):(1'h0)] reg1652 = (1'h0);
  reg [(5'h15):(1'h0)] reg1651 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1650 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1649 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1648 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1646 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1644 = (1'h0);
  reg [(4'h8):(1'h0)] reg1643 = (1'h0);
  reg [(2'h3):(1'h0)] reg1642 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1641 = (1'h0);
  reg [(4'hb):(1'h0)] reg1637 = (1'h0);
  reg [(5'h10):(1'h0)] reg1636 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1634 = (1'h0);
  reg [(3'h4):(1'h0)] reg1632 = (1'h0);
  reg [(4'hc):(1'h0)] reg1630 = (1'h0);
  reg [(5'h18):(1'h0)] reg1629 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1628 = (1'h0);
  reg [(4'h9):(1'h0)] reg1626 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1624 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1623 = (1'h0);
  reg [(2'h3):(1'h0)] reg1622 = (1'h0);
  reg [(3'h4):(1'h0)] reg1619 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1618 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1617 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1616 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1615 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1614 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1613 = (1'h0);
  reg [(4'hf):(1'h0)] reg1612 = (1'h0);
  reg [(4'hd):(1'h0)] reg1611 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1610 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar1604 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1602 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar677 = (1'h0);
  reg [(5'h14):(1'h0)] reg676 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg674 = (1'h0);
  reg [(4'hc):(1'h0)] forvar673 = (1'h0);
  reg [(5'h10):(1'h0)] forvar671 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg669 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar662 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg69 = (1'h0);
  reg [(3'h4):(1'h0)] forvar67 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg66 = (1'h0);
  reg [(5'h11):(1'h0)] reg65 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg60 = (1'h0);
  assign y = {wire1685,
                 wire1601,
                 wire1599,
                 wire659,
                 wire70,
                 wire1723,
                 wire1724,
                 wire1735,
                 reg1739,
                 reg1738,
                 reg1734,
                 reg1730,
                 reg1729,
                 reg1727,
                 reg1720,
                 reg1719,
                 reg1718,
                 reg1716,
                 reg1715,
                 reg1713,
                 reg1712,
                 reg1710,
                 reg1709,
                 reg1706,
                 reg1705,
                 reg1704,
                 reg1702,
                 reg1701,
                 reg1700,
                 reg1699,
                 reg1696,
                 reg1695,
                 reg1689,
                 reg678,
                 reg675,
                 reg672,
                 reg670,
                 reg668,
                 reg667,
                 reg666,
                 reg664,
                 reg663,
                 reg661,
                 reg68,
                 reg64,
                 reg63,
                 reg61,
                 reg59,
                 reg1603,
                 reg1605,
                 reg1606,
                 reg1607,
                 reg1608,
                 reg1609,
                 reg1620,
                 reg1621,
                 reg1625,
                 reg1627,
                 reg1631,
                 reg1633,
                 reg1635,
                 reg1638,
                 reg1639,
                 reg1640,
                 reg1645,
                 reg1647,
                 reg1654,
                 reg1656,
                 reg1657,
                 reg1658,
                 reg1659,
                 reg1664,
                 reg1665,
                 reg1666,
                 reg1670,
                 reg1672,
                 reg1674,
                 reg1676,
                 reg1684,
                 reg1737,
                 reg1733,
                 forvar1732,
                 reg1731,
                 reg1728,
                 forvar1726,
                 forvar1725,
                 reg1722,
                 reg1721,
                 reg1717,
                 reg1714,
                 reg1711,
                 reg1708,
                 reg1707,
                 reg1703,
                 reg1698,
                 forvar1697,
                 reg1690,
                 reg1697,
                 forvar1696,
                 reg1694,
                 reg1693,
                 reg1692,
                 reg1691,
                 forvar1690,
                 reg1688,
                 forvar1687,
                 reg1683,
                 reg1682,
                 reg1681,
                 reg1680,
                 reg1679,
                 reg1678,
                 reg1677,
                 reg1675,
                 reg1673,
                 reg1671,
                 reg1669,
                 reg1668,
                 reg1667,
                 reg1663,
                 reg1662,
                 reg1661,
                 reg1660,
                 reg1655,
                 reg1653,
                 reg1652,
                 reg1651,
                 reg1650,
                 reg1649,
                 reg1648,
                 forvar1646,
                 forvar1644,
                 reg1643,
                 reg1642,
                 reg1641,
                 reg1637,
                 reg1636,
                 reg1634,
                 reg1632,
                 reg1630,
                 reg1629,
                 reg1628,
                 reg1626,
                 reg1624,
                 reg1623,
                 reg1622,
                 reg1619,
                 reg1618,
                 forvar1617,
                 forvar1616,
                 reg1615,
                 reg1614,
                 forvar1613,
                 reg1612,
                 reg1611,
                 reg1610,
                 forvar1604,
                 forvar1602,
                 forvar677,
                 reg676,
                 reg674,
                 forvar673,
                 forvar671,
                 reg669,
                 reg665,
                 forvar662,
                 reg69,
                 forvar67,
                 reg66,
                 reg65,
                 reg62,
                 reg60,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire55)
        begin
          reg59 <= ($signed(((-(wire54 | wire54)) ?
              wire57 : wire55[(2'h2):(2'h2)])) > {(^~wire57[(4'ha):(3'h5)])});
          reg60 = wire58[(1'h1):(1'h1)];
          reg61 <= $signed($unsigned($unsigned(((8'ha4) ?
              $unsigned(wire54) : (^~wire58)))));
          if ($signed(wire57))
            begin
              reg62 = wire57[(3'h6):(1'h0)];
              reg63 <= reg60[(4'h8):(3'h6)];
            end
          else
            begin
              reg62 = ($signed(wire55) ?
                  (reg60 ?
                      ($unsigned(wire55[(3'h4):(1'h1)]) ^~ reg62[(2'h2):(1'h0)]) : wire56[(3'h7):(3'h4)]) : $unsigned((((reg63 ?
                          wire54 : wire57) <= (wire54 ? reg63 : (7'h44))) ?
                      wire54 : $signed(reg59))));
            end
        end
      else
        begin
          reg59 <= (($unsigned(reg59) ?
                  wire55 : {$signed(wire58[(1'h0):(1'h0)])}) ?
              (wire54 ?
                  $unsigned((8'hb5)) : (~^$unsigned((reg59 ?
                      wire57 : reg59)))) : reg60[(4'hf):(4'ha)]);
          reg61 <= (({reg62} <= wire54) ? wire56 : {$signed(wire58)});
          if ((+(reg61 - $unsigned($signed({(8'hb2)})))))
            begin
              reg63 <= (8'hae);
              reg64 <= ($signed($signed($unsigned(reg63))) ^ reg63);
              reg65 = reg62[(4'h9):(3'h6)];
            end
          else
            begin
              reg63 <= (^~wire57[(2'h3):(1'h1)]);
              reg64 <= reg63;
            end
          reg66 = (|(reg60 >> $unsigned(reg62[(4'h8):(2'h3)])));
          for (forvar67 = (1'h0); (forvar67 < (1'h0)); forvar67 = (forvar67 + (1'h1)))
            begin
              reg68 <= reg66;
              reg69 = {wire58, $signed(reg68[(1'h0):(1'h0)])};
            end
        end
    end
  assign wire70 = $unsigned(($signed(wire58) == (((!reg68) >> $signed((8'ha1))) != (+(wire54 && (8'hbe))))));
  module71 #() modinst660 (.clk(clk), .y(wire659), .wire75(wire70), .wire73(wire58), .wire72(reg68), .wire74(reg63));
  always
    @(posedge clk) begin
      reg661 <= $signed((|$signed($signed($signed(reg59)))));
      for (forvar662 = (1'h0); (forvar662 < (1'h1)); forvar662 = (forvar662 + (1'h1)))
        begin
          if (reg68[(3'h7):(1'h1)])
            begin
              reg663 <= $unsigned($signed((^~(+(~^wire54)))));
              reg664 <= wire57[(4'h8):(2'h3)];
              reg665 = $signed((~|wire55[(4'he):(3'h7)]));
            end
          else
            begin
              reg665 = $unsigned(($unsigned(((wire57 ? wire57 : reg61) ?
                  reg59[(1'h0):(1'h0)] : ((8'hbb) ?
                      reg63 : (8'hae)))) <<< $signed(wire57[(4'ha):(4'h9)])));
              reg666 <= (($unsigned({reg63[(2'h2):(1'h0)]}) ?
                      ($signed(((8'ha4) >> reg664)) ?
                          reg665[(5'h12):(5'h12)] : {{wire659, reg661},
                              ((7'h46) || wire55)}) : ($unsigned($unsigned(reg61)) ?
                          $signed(reg661) : $unsigned($signed(reg68)))) ?
                  $unsigned(reg59) : reg63[(2'h3):(2'h2)]);
              reg667 <= {reg61, $unsigned(reg68)};
              reg668 <= (8'hbc);
              reg669 = $unsigned(reg663[(4'hd):(3'h4)]);
            end
          reg670 <= $signed((8'haf));
          for (forvar671 = (1'h0); (forvar671 < (3'h4)); forvar671 = (forvar671 + (1'h1)))
            begin
              reg672 <= (^~{$unsigned({$unsigned(reg59)})});
            end
          for (forvar673 = (1'h0); (forvar673 < (1'h0)); forvar673 = (forvar673 + (1'h1)))
            begin
              reg674 = reg68;
              reg675 <= $unsigned(({$signed(wire56)} ~^ $unsigned((~(~wire57)))));
              reg676 = (|{($unsigned((reg672 ? forvar662 : reg675)) ?
                      ((reg664 ? (8'h9f) : reg669) ?
                          (reg674 ^ reg666) : $unsigned(wire57)) : $signed((wire54 ?
                          reg670 : reg672)))});
            end
          for (forvar677 = (1'h0); (forvar677 < (2'h2)); forvar677 = (forvar677 + (1'h1)))
            begin
              reg678 <= forvar662[(4'he):(4'hb)];
            end
        end
    end
  module679 #() modinst1600 (.clk(clk), .wire683(reg668), .y(wire1599), .wire684(reg59), .wire681(reg675), .wire680(reg64), .wire682(reg68));
  assign wire1601 = (reg661 && reg672[(4'h9):(4'h9)]);
  always
    @(posedge clk) begin
      for (forvar1602 = (1'h0); (forvar1602 < (2'h3)); forvar1602 = (forvar1602 + (1'h1)))
        begin
          reg1603 <= ((reg61[(2'h2):(2'h2)] ?
              ((|$unsigned(reg59)) ^~ forvar1602[(4'h9):(4'h9)]) : {$signed($unsigned(reg64)),
                  $unsigned(reg68)}) * $unsigned($signed($unsigned((wire1599 - reg675)))));
          for (forvar1604 = (1'h0); (forvar1604 < (1'h1)); forvar1604 = (forvar1604 + (1'h1)))
            begin
              reg1605 <= (&(^~$unsigned(reg667[(2'h2):(1'h1)])));
              reg1606 <= (reg661 > {forvar1604, (|wire57)});
              reg1607 <= {(($unsigned((|reg672)) ?
                          $signed(forvar1604) : reg678[(3'h4):(1'h0)]) ?
                      wire70[(5'h11):(1'h1)] : reg68[(5'h12):(3'h7)])};
              reg1608 <= $unsigned(({$signed(wire659[(2'h3):(1'h1)])} ?
                  ((wire56 ?
                          (reg1603 ? wire1599 : (8'ha3)) : (reg668 >> reg64)) ?
                      ((~(8'hb9)) ?
                          wire56[(3'h6):(3'h5)] : $signed(wire70)) : ((8'hbc) ?
                          (reg664 ~^ wire57) : $unsigned(reg59))) : reg661[(5'h10):(4'hf)]));
            end
          if ($signed($unsigned((reg670[(5'h10):(4'he)] ?
              ((&reg1603) ?
                  (reg678 ? reg1606 : (8'hbd)) : (8'hb5)) : (!(7'h44))))))
            begin
              reg1609 <= $unsigned($signed(((!(reg667 <= reg667)) ?
                  wire1601 : $unsigned(reg1607))));
              reg1610 = forvar1602[(3'h5):(3'h5)];
              reg1611 = {reg1605};
              reg1612 = (~^reg664[(3'h7):(3'h7)]);
            end
          else
            begin
              reg1610 = wire1601;
            end
          for (forvar1613 = (1'h0); (forvar1613 < (2'h2)); forvar1613 = (forvar1613 + (1'h1)))
            begin
              reg1614 = $unsigned(($signed(reg1610[(2'h2):(2'h2)]) ?
                  reg1605[(2'h2):(2'h2)] : wire659[(2'h2):(1'h0)]));
              reg1615 = (((~&{$unsigned(reg1612)}) - wire659[(3'h5):(3'h5)]) || (reg1606[(1'h0):(1'h0)] > ((^$signed(wire56)) - {reg61,
                  (|reg68)})));
            end
        end
      for (forvar1616 = (1'h0); (forvar1616 < (1'h0)); forvar1616 = (forvar1616 + (1'h1)))
        begin
          for (forvar1617 = (1'h0); (forvar1617 < (2'h2)); forvar1617 = (forvar1617 + (1'h1)))
            begin
              reg1618 = {reg63,
                  $signed((forvar1617[(3'h4):(2'h2)] ?
                      $unsigned((forvar1617 ? reg1612 : (7'h44))) : reg670))};
              reg1619 = reg1606;
            end
          reg1620 <= $signed(forvar1616);
          if (reg1603)
            begin
              reg1621 <= ($signed((((7'h46) ?
                      (reg1611 ?
                          reg1606 : reg1608) : ((7'h41) & wire54)) + reg1615)) ?
                  $unsigned($unsigned(($signed(reg1615) && $unsigned(reg1612)))) : (($unsigned({(8'h9c),
                          wire58}) ^~ $unsigned(wire54[(2'h3):(1'h0)])) ?
                      $unsigned(((~forvar1613) <<< (reg1607 ?
                          wire659 : wire1599))) : (reg1603 ?
                          {$unsigned(forvar1616)} : $signed(forvar1617))));
              reg1622 = (^(+reg1610[(1'h0):(1'h0)]));
              reg1623 = {$signed((^~(~(reg1610 ? (8'hac) : reg1614)))),
                  wire659};
              reg1624 = $unsigned({forvar1617[(4'hd):(3'h6)]});
            end
          else
            begin
              reg1621 <= wire659[(4'hd):(3'h4)];
              reg1625 <= $signed($unsigned({(~(reg1610 <= reg1619))}));
              reg1626 = $unsigned({((reg1623[(1'h0):(1'h0)] ?
                          $signed(wire659) : $signed((8'h9e))) ?
                      (+forvar1602[(3'h5):(3'h5)]) : (8'hae))});
              reg1627 <= $signed($unsigned((wire659 + reg1603[(2'h3):(1'h1)])));
              reg1628 = ((((reg59[(2'h2):(1'h1)] >= reg1620) ?
                      ((&forvar1602) ^ (reg663 < (7'h46))) : {$signed(wire57),
                          reg63[(3'h4):(2'h2)]}) != $unsigned(((reg666 ?
                          reg1611 : reg663) ?
                      reg1607 : $signed((8'had))))) ?
                  $signed((|$unsigned($signed(reg1611)))) : (~|forvar1617));
            end
        end
      if (({reg1614[(2'h3):(1'h0)], ((|$signed(reg1625)) > reg1627)} ?
          ($signed((reg1625 * $signed(wire659))) ?
              $signed((~&$signed((8'hb7)))) : ($signed({(7'h46), reg1619}) ?
                  $signed((reg64 ^~ reg1627)) : $signed($signed((8'hbe))))) : reg1612[(4'h8):(1'h1)]))
        begin
          if (reg1620[(4'h8):(1'h1)])
            begin
              reg1629 = (+reg1623);
              reg1630 = $signed($signed(reg1622));
              reg1631 <= $unsigned($unsigned(($unsigned((+wire1599)) ?
                  $unsigned(((8'ha2) < reg1623)) : (reg1626[(3'h4):(1'h0)] <= {reg675}))));
              reg1632 = $unsigned(((reg1629 >>> reg1610) ^~ $signed($signed((reg670 > (8'ha8))))));
              reg1633 <= ($signed($unsigned($unsigned(reg1621[(4'hc):(4'h9)]))) ?
                  reg1624 : (reg675[(3'h6):(2'h2)] ?
                      ($unsigned(wire56) * $unsigned($unsigned(reg1620))) : {(|reg1632[(3'h4):(3'h4)])}));
            end
          else
            begin
              reg1629 = reg1627[(1'h0):(1'h0)];
              reg1630 = (($signed($unsigned((~forvar1613))) ?
                  $signed(reg1627[(1'h1):(1'h1)]) : reg1624) | ((reg59[(3'h6):(3'h5)] & $signed((-(8'haf)))) + {$unsigned(((8'hae) >= reg1630)),
                  $signed($signed(reg663))}));
              reg1631 <= {wire1599,
                  ((+reg1605) ?
                      {$signed((reg1611 || reg1605)),
                          (8'h9c)} : reg667[(4'hc):(1'h1)])};
              reg1633 <= $signed(reg1603);
            end
        end
      else
        begin
          if ((8'hbe))
            begin
              reg1631 <= reg59[(3'h7):(3'h5)];
              reg1632 = $unsigned((((-(reg59 ? reg1631 : wire55)) ?
                      $signed(reg1605) : (8'ha1)) ?
                  forvar1604 : (((forvar1602 ? reg1630 : reg1633) ?
                          (reg1623 - (8'hb7)) : reg675) ?
                      {$signed(reg64)} : ({reg1614} >> reg1630[(4'h9):(3'h4)]))));
              reg1633 <= wire1599;
              reg1634 = $unsigned((8'hb6));
              reg1635 <= $signed((!(reg661 || $signed({reg675}))));
            end
          else
            begin
              reg1631 <= wire70;
              reg1632 = $signed(reg667);
              reg1634 = (((((!wire55) ?
                              $signed(forvar1613) : $unsigned(reg678)) ?
                          {reg1631,
                              (reg68 ?
                                  reg667 : reg666)} : reg666[(5'h14):(5'h14)]) ?
                      {((reg1632 ? (8'hb9) : reg1635) ? (8'hb7) : (7'h48)),
                          (~|$unsigned(reg1626))} : reg664) ?
                  (+reg666) : (~reg664[(4'h9):(1'h0)]));
              reg1635 <= $unsigned($unsigned(reg59));
            end
          if (($signed((((&reg1622) | $unsigned(reg661)) ?
              ((reg1627 ? reg1624 : reg1606) >>> reg1618) : ((reg61 ?
                  (8'hb7) : reg672) ^~ (-(8'hb3))))) || {((~&{reg666,
                      reg1623}) ?
                  ($unsigned(reg1620) + $unsigned(reg1607)) : (|$unsigned(reg1635)))}))
            begin
              reg1636 = $unsigned((wire55[(4'ha):(1'h1)] ?
                  $signed(((reg68 ? (8'h9f) : wire1599) ?
                      (reg1619 ? forvar1602 : reg1629) : {reg1619})) : wire58));
              reg1637 = ($signed((((8'hab) ?
                  reg1605 : $unsigned(reg1608)) & $unsigned(reg1623))) && (+(({wire58} ?
                  reg1606[(3'h5):(2'h2)] : $unsigned(wire659)) ^ reg1615[(3'h5):(2'h3)])));
              reg1638 <= $unsigned($signed($unsigned(forvar1604[(2'h3):(1'h1)])));
              reg1639 <= ((($signed($signed(reg1622)) ?
                      $signed({reg59,
                          wire56}) : (wire1599[(3'h4):(1'h0)] || $signed(wire58))) ?
                  (reg1603 ?
                      reg664[(2'h2):(2'h2)] : (~^(&reg64))) : reg1625[(3'h5):(1'h1)]) >>> $unsigned($signed(({forvar1613} + $unsigned(wire58)))));
              reg1640 <= $signed(forvar1617[(4'hd):(4'hb)]);
            end
          else
            begin
              reg1636 = {reg1623,
                  ((&$signed(reg661)) ?
                      {{$signed(forvar1604),
                              (reg1614 < reg1621)}} : (reg668 << forvar1613))};
              reg1638 <= ($unsigned($signed(reg1633)) ?
                  {{((^~reg1638) <= (^~(8'ha9))), reg1619},
                      ($unsigned(reg1614[(2'h2):(1'h1)]) >> reg63[(3'h5):(3'h5)])} : $signed((~|((reg672 ?
                      reg666 : (7'h44)) == reg1606))));
            end
          if (reg1603)
            begin
              reg1641 = ($signed((8'hae)) != (reg1612[(4'ha):(1'h0)] ?
                  $signed(((reg668 ~^ wire55) && $signed(reg1606))) : $unsigned($unsigned((reg1637 ?
                      forvar1604 : wire55)))));
              reg1642 = reg1629[(5'h17):(5'h10)];
            end
          else
            begin
              reg1641 = $unsigned((forvar1604 ?
                  reg1640[(1'h1):(1'h0)] : $unsigned((~&(~^wire54)))));
              reg1642 = $signed((($signed((7'h4a)) & reg1632) <= wire56));
            end
          reg1643 = reg63[(3'h6):(2'h3)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar1644 = (1'h0); (forvar1644 < (2'h3)); forvar1644 = (forvar1644 + (1'h1)))
        begin
          reg1645 <= wire1599;
          for (forvar1646 = (1'h0); (forvar1646 < (2'h2)); forvar1646 = (forvar1646 + (1'h1)))
            begin
              reg1647 <= (^(!$unsigned(({reg670} ?
                  $signed(reg1631) : (wire56 <= wire659)))));
              reg1648 = (~^(|{wire58[(5'h12):(4'h8)]}));
              reg1649 = (-((((8'hb7) ^~ {reg1607,
                      reg678}) > reg1627[(1'h1):(1'h0)]) ?
                  (8'had) : reg59[(3'h6):(3'h6)]));
              reg1650 = $signed($signed((((^~reg675) > (reg1603 ?
                  reg1608 : reg667)) < $signed(reg667[(4'hf):(3'h4)]))));
              reg1651 = (~^reg1631);
            end
          if ($signed($signed(((reg1606[(1'h0):(1'h0)] ~^ ((8'ha8) ?
              reg668 : reg664)) <= wire1599))))
            begin
              reg1652 = reg1607;
              reg1653 = ($unsigned($unsigned(($unsigned((8'ha3)) ?
                      reg1649[(3'h7):(2'h2)] : reg1652))) ?
                  wire1599 : $signed($unsigned(reg667[(2'h2):(1'h1)])));
            end
          else
            begin
              reg1654 <= ($unsigned((($unsigned(reg1605) ? reg670 : (+wire57)) ?
                  {{(8'hb0)}} : reg1645[(4'ha):(4'ha)])) << (^reg661));
              reg1655 = $signed($signed($signed((~&$unsigned(reg63)))));
              reg1656 <= (reg1651 >> reg1633);
              reg1657 <= (reg670 ?
                  (reg1620 ?
                      $unsigned(($signed(reg1640) ?
                          (&wire55) : (&wire55))) : reg1639[(4'hc):(2'h2)]) : reg678);
              reg1658 <= ({$signed({(wire57 > forvar1644),
                      $unsigned(wire1601)}),
                  reg1651} <= {reg672[(4'hc):(3'h7)], wire57});
            end
          if ({(((reg1652 ?
                  (reg1606 ? reg1631 : reg1621) : (reg1658 ?
                      reg675 : reg1649)) & (^~(~|reg1651))) >= (^~reg1609[(2'h3):(1'h1)])),
              {$unsigned($signed($signed((8'hac)))),
                  (~^(reg1631 <<< $unsigned(wire56)))}})
            begin
              reg1659 <= $unsigned(reg668[(5'h13):(2'h3)]);
            end
          else
            begin
              reg1660 = ($signed(wire70) <<< (^~reg63[(2'h2):(1'h0)]));
              reg1661 = (~|{$signed((~^(reg1609 ? reg1648 : (8'hbb)))),
                  {$unsigned(wire56[(3'h6):(2'h3)]), reg1656[(1'h0):(1'h0)]}});
              reg1662 = (&(reg1631 >>> wire70[(5'h13):(5'h11)]));
              reg1663 = $signed((!(!$unsigned((~^forvar1646)))));
              reg1664 <= (^~reg1647);
            end
        end
      reg1665 <= (($signed((reg1655[(4'h9):(3'h4)] ?
                  $unsigned(reg1633) : $unsigned(reg1608))) ?
              $unsigned({$signed(reg1608),
                  $unsigned(reg1650)}) : wire54[(4'hd):(3'h7)]) ?
          reg675 : (wire58 ?
              reg1603[(3'h4):(1'h0)] : ($unsigned((reg663 ?
                  reg1609 : reg661)) - $unsigned((reg1631 >>> reg678)))));
    end
  always
    @(posedge clk) begin
      reg1666 <= $signed((reg666 == (reg1638 * ((^~reg1656) & $unsigned(reg1605)))));
      reg1667 = reg1640;
      reg1668 = $signed(reg1667);
      if (reg1638[(1'h0):(1'h0)])
        begin
          reg1669 = $signed(wire1601);
        end
      else
        begin
          reg1670 <= $unsigned(((~$signed(((8'hbc) ? reg1627 : reg1667))) ?
              $unsigned($unsigned(reg672)) : (({reg1667} || $signed((8'had))) >= reg1638)));
          reg1671 = $unsigned(reg661);
          if (((reg1647 ?
                  (+{(wire58 ^~ (7'h40)),
                      (reg666 || reg664)}) : ($unsigned((reg64 ?
                      reg666 : (8'hb2))) >= (~^((8'hb6) ? wire58 : wire56)))) ?
              $unsigned(($unsigned(reg1668[(2'h2):(2'h2)]) ?
                  reg1654 : $unsigned((~^reg1633)))) : $unsigned($signed({$signed(reg1627)}))))
            begin
              reg1672 <= {$unsigned({wire659[(2'h3):(2'h3)],
                      ((reg1635 * reg1621) ? $unsigned((8'hb3)) : reg1666)}),
                  reg678};
              reg1673 = (~|($unsigned($unsigned($signed(wire57))) ?
                  reg1635[(3'h5):(2'h2)] : {((^~(7'h41)) ?
                          reg1666 : (~^(8'ha6))),
                      ($signed(reg666) ?
                          $unsigned(wire1599) : (reg1635 ~^ reg1668))}));
            end
          else
            begin
              reg1672 <= reg64[(4'hf):(3'h6)];
              reg1674 <= (^~$unsigned(($unsigned((~^reg675)) <= $signed((~(8'ha0))))));
            end
          if (({(~&{$unsigned(reg1664)})} >= reg1603))
            begin
              reg1675 = ($signed(reg1621) ?
                  ($unsigned(($signed(reg1621) ?
                          $signed(reg678) : (reg1640 > reg1668))) ?
                      $signed($signed(wire1599)) : $signed(reg1665[(5'h12):(3'h4)])) : reg1659[(3'h6):(2'h2)]);
              reg1676 <= ($unsigned(({reg1605} ?
                  (wire659 ?
                      reg61[(2'h3):(1'h0)] : reg1667) : (~|$signed(reg664)))) >= $signed(((~reg1620) && wire57[(2'h3):(1'h0)])));
              reg1677 = ((reg1625 ?
                      $unsigned(reg1657[(3'h4):(1'h1)]) : (!$unsigned(reg1659[(4'ha):(3'h7)]))) ?
                  $unsigned((8'h9d)) : ($signed((8'hb2)) ?
                      ({((8'hb7) ?
                              reg1674 : reg59)} <<< reg1608[(5'h10):(4'hc)]) : ($unsigned(reg1603[(3'h5):(1'h1)]) ?
                          $signed((wire56 ? wire1599 : reg63)) : reg670)));
              reg1678 = ({(7'h45)} ?
                  (((reg1638 ? (reg63 ? reg1677 : reg678) : (+reg1635)) ?
                          $signed($signed(reg1608)) : (~^$unsigned(wire57))) ?
                      (~|reg1676) : $unsigned({(7'h4a)})) : {((reg1607 >= $unsigned(reg1654)) ?
                          (&(^reg1656)) : $signed(reg1677))});
            end
          else
            begin
              reg1676 <= reg1609;
              reg1677 = ({$unsigned(((^~wire54) ?
                      (reg1667 ?
                          reg68 : reg663) : wire70[(5'h14):(4'hd)]))} ^ reg1678[(1'h0):(1'h0)]);
              reg1678 = (8'hb5);
              reg1679 = {reg678[(4'h8):(1'h0)], reg61[(1'h1):(1'h1)]};
            end
          reg1680 = (reg1671 ? reg1654 : reg1633);
        end
    end
  always
    @(posedge clk) begin
      reg1681 = reg1605;
      reg1682 = (8'ha9);
      reg1683 = ($unsigned({({reg1654} ?
              $signed(reg1638) : (reg672 - reg678))}) ^ ((+reg678[(3'h7):(3'h6)]) ?
          ({$signed(reg1607), $unsigned(reg1657)} ?
              (7'h46) : ($unsigned(reg668) ?
                  $unsigned(reg1659) : $unsigned(reg1674))) : reg672[(5'h10):(2'h3)]));
      reg1684 <= (((reg1603 ?
              wire1599[(3'h4):(1'h1)] : ($unsigned(reg1603) ?
                  $unsigned(reg1654) : $signed(reg672))) >> reg1681) ?
          $signed(((8'h9c) ?
              (^{reg1657}) : (reg1666 ?
                  reg667 : ((8'h9d) >>> reg64)))) : $signed($signed($signed((|reg672)))));
    end
  module195 #() modinst1686 (.wire196(reg661), .y(wire1685), .wire197(wire55), .clk(clk), .wire199(reg668), .wire198(reg1672));
  always
    @(posedge clk) begin
      for (forvar1687 = (1'h0); (forvar1687 < (2'h2)); forvar1687 = (forvar1687 + (1'h1)))
        begin
          reg1688 = (~|$signed(($unsigned((reg1665 ? reg1603 : reg666)) ?
              (reg675 <<< reg1635[(2'h3):(2'h2)]) : $signed(wire1599))));
        end
      if (reg668)
        begin
          reg1689 <= {reg1654[(1'h0):(1'h0)]};
          for (forvar1690 = (1'h0); (forvar1690 < (1'h1)); forvar1690 = (forvar1690 + (1'h1)))
            begin
              reg1691 = wire70;
              reg1692 = forvar1690;
              reg1693 = (!wire54[(4'he):(1'h1)]);
              reg1694 = ($unsigned(($unsigned(wire70[(5'h12):(3'h5)]) ?
                      ($unsigned(reg1665) ?
                          (reg1656 >>> reg1608) : reg1621) : wire1599[(3'h4):(2'h3)])) ?
                  $signed(((^~reg1647[(3'h6):(3'h5)]) ?
                      $unsigned($signed(reg678)) : reg672)) : (((|((8'ha3) ?
                      reg63 : reg1635)) <<< $signed($signed(wire1685))) | ({(reg672 >= reg1625)} & {(wire1601 >> wire1685),
                      ((8'hb7) == reg1638)})));
              reg1695 <= (^~reg1609[(5'h10):(4'ha)]);
            end
          for (forvar1696 = (1'h0); (forvar1696 < (1'h0)); forvar1696 = (forvar1696 + (1'h1)))
            begin
              reg1697 = (&$signed(reg1670[(2'h2):(2'h2)]));
            end
        end
      else
        begin
          if (($unsigned(reg663[(2'h2):(1'h1)]) ?
              reg1645 : (~|reg1691[(4'hc):(1'h1)])))
            begin
              reg1689 <= ($signed(reg68[(1'h1):(1'h0)]) != (~|(reg1659 != $unsigned($unsigned(reg1664)))));
              reg1690 = ((~^((~&(reg1676 ~^ reg675)) ?
                      ($signed(reg1654) && $unsigned(reg1684)) : $signed((~^reg1670)))) ?
                  (reg1609 ?
                      ($signed((reg1657 ~^ (8'hac))) > ((reg1639 ?
                          reg68 : reg1608) && $signed(reg1645))) : reg1694) : reg661);
            end
          else
            begin
              reg1690 = (({$signed((!reg1665)),
                          (reg1606[(3'h7):(3'h5)] == $unsigned(reg1625))} ?
                      reg1690 : $signed($unsigned(reg1664))) ?
                  (((!$signed(reg1621)) >= (^(reg668 ?
                      wire1685 : reg1605))) >= wire1685) : reg1684[(1'h1):(1'h1)]);
              reg1695 <= (wire659 ^~ $unsigned((((~^reg1621) ?
                  reg1631 : $unsigned((8'ha6))) - reg1697)));
              reg1696 <= $unsigned($signed($signed(reg1676[(4'h8):(2'h3)])));
            end
          for (forvar1697 = (1'h0); (forvar1697 < (1'h0)); forvar1697 = (forvar1697 + (1'h1)))
            begin
              reg1698 = wire1599[(3'h4):(2'h2)];
              reg1699 <= ($signed((^~(reg1657 ?
                  (reg1645 ?
                      wire659 : (8'h9c)) : (^~reg1656)))) != $signed({reg1693[(2'h2):(2'h2)]}));
              reg1700 <= $signed(reg1657);
              reg1701 <= $unsigned(reg68[(5'h13):(5'h10)]);
              reg1702 <= {(reg1676[(3'h6):(1'h0)] ?
                      $unsigned($signed(reg1605[(1'h0):(1'h0)])) : ($signed(reg678[(3'h4):(1'h0)]) >>> $unsigned(wire1685[(4'h9):(3'h6)]))),
                  reg61};
            end
        end
      if ((^~$signed($signed($signed(wire55)))))
        begin
          if ((reg1694 + $signed((~|(reg1625 >> reg1698[(4'hf):(3'h6)])))))
            begin
              reg1703 = (8'h9c);
            end
          else
            begin
              reg1704 <= (-reg1699[(4'hd):(3'h6)]);
              reg1705 <= $signed(((~|(!wire54)) * wire57));
              reg1706 <= reg1666[(1'h1):(1'h1)];
            end
          if ({(^($signed(reg1705[(3'h6):(2'h2)]) ^ (&(reg1639 ?
                  reg1609 : reg68)))),
              reg670[(5'h12):(5'h12)]})
            begin
              reg1707 = $unsigned(($signed(($unsigned(reg1700) ?
                      (-reg1664) : reg1700)) ?
                  $signed($unsigned((reg1607 ?
                      wire58 : reg1692))) : $signed((~|reg1645[(4'hb):(4'h9)]))));
              reg1708 = $signed($unsigned((!$unsigned(wire1685))));
              reg1709 <= $signed($signed((^~$signed(reg661[(4'h8):(3'h4)]))));
              reg1710 <= reg1694;
            end
          else
            begin
              reg1709 <= $unsigned((-{(!forvar1696[(2'h2):(1'h1)])}));
              reg1710 <= reg1620[(2'h2):(2'h2)];
            end
          if (($unsigned({reg1666[(3'h7):(2'h2)],
              $unsigned(forvar1696)}) & reg1664))
            begin
              reg1711 = (reg1607[(2'h2):(2'h2)] ?
                  reg1656[(3'h5):(2'h2)] : $unsigned((((reg59 ?
                      forvar1697 : reg1704) == (+reg1691)) >> $unsigned($unsigned(reg672)))));
            end
          else
            begin
              reg1711 = (($signed(((reg63 + reg1674) ?
                          $unsigned((8'hb3)) : ((8'ha5) & wire57))) ?
                      reg1659 : $signed(wire659[(3'h5):(2'h2)])) ?
                  reg1692[(3'h4):(3'h4)] : $signed($unsigned({$unsigned(reg668)})));
              reg1712 <= reg675[(2'h3):(1'h1)];
              reg1713 <= (8'ha7);
              reg1714 = (reg670 ?
                  {(~$unsigned((reg1605 <<< reg672))),
                      ({$signed(reg1698)} ?
                          ($unsigned(reg1712) ?
                              {reg1640,
                                  reg1656} : reg1609[(4'he):(3'h7)]) : (~$signed(reg1690)))} : (wire56[(3'h6):(2'h3)] ?
                      reg1665 : $signed($unsigned((wire70 ?
                          reg1666 : reg68)))));
            end
          reg1715 <= {($unsigned(((reg1672 ? (8'ha9) : (8'hac)) ~^ (reg678 ?
                      reg68 : reg1647))) ?
                  reg1666[(4'hb):(1'h1)] : $unsigned(((reg1633 ?
                      reg1654 : forvar1690) || (reg672 || reg1640))))};
          reg1716 <= (reg1621 ?
              $signed(($unsigned((!reg1672)) ^~ (~|reg61))) : $signed($unsigned((&(8'h9c)))));
        end
      else
        begin
          reg1703 = ($signed((8'ha6)) ?
              (-{wire58}) : $unsigned((reg667 ? (8'hae) : reg1702)));
          if (wire1601[(2'h2):(1'h0)])
            begin
              reg1707 = $signed($signed(reg1714));
              reg1708 = ((&$unsigned(((!reg666) ?
                      $unsigned(reg1674) : (reg1620 ? (7'h44) : reg1709)))) ?
                  ({reg1664} ?
                      reg1672 : {$unsigned(reg63[(1'h1):(1'h1)]),
                          ((8'haa) >> reg1672[(4'hb):(1'h0)])}) : ($unsigned((reg1713[(1'h1):(1'h1)] << $unsigned(reg1656))) ?
                      $signed($signed($unsigned(reg1707))) : $signed($signed($unsigned(reg1712)))));
              reg1711 = $unsigned($unsigned($signed(reg666[(1'h1):(1'h0)])));
              reg1712 <= (^$signed(reg68));
            end
          else
            begin
              reg1704 <= (^reg1640[(3'h4):(2'h3)]);
              reg1705 <= (&{((|wire1685[(4'hb):(3'h5)]) ?
                      $unsigned(reg1645[(4'hc):(1'h0)]) : ($signed(reg1714) * reg663[(4'h9):(2'h2)])),
                  (reg1664[(4'h8):(2'h3)] & $unsigned(reg675))});
              reg1707 = $unsigned(wire55[(4'he):(4'ha)]);
              reg1709 <= (+reg1620);
            end
          reg1714 = $signed($unsigned($signed(wire57[(3'h7):(3'h6)])));
          if ((reg678 != reg1688))
            begin
              reg1715 <= (7'h40);
              reg1716 <= (~|$unsigned(reg1706[(1'h0):(1'h0)]));
              reg1717 = $unsigned($unsigned((reg1712 ?
                  reg1694[(3'h7):(3'h6)] : $signed($signed(reg1700)))));
            end
          else
            begin
              reg1717 = reg678;
              reg1718 <= (^({((reg1716 && reg1645) ?
                      $unsigned(reg1688) : (reg1645 >> (7'h47)))} | (+($signed((8'hae)) ?
                  $unsigned((8'haa)) : reg1715))));
              reg1719 <= $signed(($signed(reg1627[(1'h0):(1'h0)]) ?
                  reg1640 : (8'haa)));
              reg1720 <= (!($signed(($unsigned(wire1599) == $signed(reg1676))) ?
                  ((((8'hb9) <= reg63) ? (+reg1691) : $signed(reg666)) ?
                      $signed((8'h9c)) : $unsigned($unsigned(reg1698))) : reg1639[(4'hc):(3'h5)]));
              reg1721 = (((^reg1647[(3'h6):(1'h1)]) ?
                      $signed((8'ha2)) : (wire70 & (-reg1638[(2'h2):(1'h1)]))) ?
                  $signed($signed(wire659[(1'h1):(1'h0)])) : reg1700[(4'h9):(3'h4)]);
            end
        end
      reg1722 = $signed(reg1645[(2'h3):(2'h3)]);
    end
  assign wire1723 = reg1670;
  assign wire1724 = $unsigned(reg678[(1'h0):(1'h0)]);
  always
    @(posedge clk) begin
      for (forvar1725 = (1'h0); (forvar1725 < (2'h2)); forvar1725 = (forvar1725 + (1'h1)))
        begin
          for (forvar1726 = (1'h0); (forvar1726 < (2'h2)); forvar1726 = (forvar1726 + (1'h1)))
            begin
              reg1727 <= reg1656[(3'h6):(3'h5)];
              reg1728 = reg1705[(4'h8):(4'h8)];
              reg1729 <= reg1639[(1'h0):(1'h0)];
              reg1730 <= $unsigned(reg1645);
              reg1731 = {(|$signed($signed($unsigned((8'ha4))))),
                  ((+reg666) == $unsigned(($unsigned(reg1638) ?
                      ((8'ha4) ? reg1670 : reg1729) : (|reg1700))))};
            end
          for (forvar1732 = (1'h0); (forvar1732 < (2'h2)); forvar1732 = (forvar1732 + (1'h1)))
            begin
              reg1733 = $unsigned({(~&$signed(reg1689)), reg1712});
            end
        end
      reg1734 <= $signed(reg1639[(4'h8):(2'h3)]);
    end
  module522 #() modinst1736 (.wire525(reg1727), .clk(clk), .wire523(reg59), .wire527(wire1685), .wire526(reg1713), .y(wire1735), .wire524(reg1658));
  always
    @(posedge clk) begin
      reg1737 = ((($signed(wire70) ?
          (8'hac) : $signed(reg1676[(4'hb):(1'h1)])) - reg1729) != wire1601[(1'h1):(1'h1)]);
      reg1738 <= (reg1639[(3'h4):(1'h1)] ?
          ($signed($signed($unsigned(reg1734))) ?
              reg1729 : reg1727) : (reg1704 ?
              $unsigned(wire70[(4'hf):(3'h5)]) : $unsigned(($signed(wire57) < (!reg670)))));
      reg1739 <= {(&(^~$signed($signed(reg1705))))};
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module679
#(parameter param1597 = (((^(((8'hbd) ? (8'h9c) : (7'h48)) >> ((7'h45) && (8'h9e)))) >= ({(^~(8'hb3))} + (^~((8'hac) >> (8'h9d))))) ? (8'ha4) : ((^~((~^(8'ha6)) ^ ((7'h42) & (8'ha3)))) && (~^(((8'h9f) ^ (8'hbf)) != ((7'h4a) ? (8'hae) : (7'h45)))))), 
parameter param1598 = (^param1597))
(y, clk, wire680, wire681, wire682, wire683, wire684);
  output wire [(32'hd51):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire680;
  input wire signed [(4'ha):(1'h0)] wire681;
  input wire signed [(4'hf):(1'h0)] wire682;
  input wire signed [(5'h13):(1'h0)] wire683;
  input wire signed [(5'h13):(1'h0)] wire684;
  wire signed [(5'h14):(1'h0)] wire1595;
  wire [(5'h14):(1'h0)] wire1593;
  wire [(3'h5):(1'h0)] wire1431;
  wire signed [(4'h9):(1'h0)] wire1337;
  wire signed [(5'h15):(1'h0)] wire1335;
  wire signed [(5'h17):(1'h0)] wire1138;
  wire signed [(3'h5):(1'h0)] wire872;
  reg [(2'h3):(1'h0)] reg1596 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1430 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1429 = (1'h0);
  reg [(4'hf):(1'h0)] reg1428 = (1'h0);
  reg [(4'hb):(1'h0)] reg1427 = (1'h0);
  reg [(5'h16):(1'h0)] reg1426 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1424 = (1'h0);
  reg [(3'h7):(1'h0)] reg1422 = (1'h0);
  reg [(5'h17):(1'h0)] reg1421 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1414 = (1'h0);
  reg [(2'h3):(1'h0)] reg1418 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1417 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1416 = (1'h0);
  reg [(5'h14):(1'h0)] reg1415 = (1'h0);
  reg [(5'h12):(1'h0)] reg1413 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1400 = (1'h0);
  reg [(4'hd):(1'h0)] reg1396 = (1'h0);
  reg [(4'he):(1'h0)] reg1412 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1408 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1407 = (1'h0);
  reg [(4'h8):(1'h0)] reg1405 = (1'h0);
  reg [(5'h10):(1'h0)] reg1402 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1401 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1398 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1397 = (1'h0);
  reg [(3'h5):(1'h0)] reg1394 = (1'h0);
  reg [(3'h6):(1'h0)] reg1393 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1392 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1390 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1388 = (1'h0);
  reg [(5'h16):(1'h0)] reg1386 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1381 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1380 = (1'h0);
  reg [(4'h9):(1'h0)] reg1376 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1374 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1373 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1371 = (1'h0);
  reg [(5'h14):(1'h0)] reg1370 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1368 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1365 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1364 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1363 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1362 = (1'h0);
  reg [(2'h3):(1'h0)] reg1361 = (1'h0);
  reg [(4'hf):(1'h0)] reg1358 = (1'h0);
  reg [(2'h3):(1'h0)] reg1355 = (1'h0);
  reg [(4'hd):(1'h0)] reg1353 = (1'h0);
  reg [(5'h17):(1'h0)] reg1351 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1350 = (1'h0);
  reg [(4'hd):(1'h0)] reg1349 = (1'h0);
  reg [(3'h6):(1'h0)] reg1345 = (1'h0);
  reg [(3'h6):(1'h0)] reg1338 = (1'h0);
  reg [(3'h4):(1'h0)] reg686 = (1'h0);
  reg [(5'h14):(1'h0)] reg688 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg691 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg693 = (1'h0);
  reg [(4'hc):(1'h0)] reg694 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg696 = (1'h0);
  reg [(4'ha):(1'h0)] reg697 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg701 = (1'h0);
  reg [(5'h11):(1'h0)] reg702 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg703 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg704 = (1'h0);
  reg signed [(4'he):(1'h0)] reg708 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg707 = (1'h0);
  reg [(5'h12):(1'h0)] reg712 = (1'h0);
  reg [(2'h3):(1'h0)] reg715 = (1'h0);
  reg signed [(4'he):(1'h0)] reg718 = (1'h0);
  reg [(5'h12):(1'h0)] reg721 = (1'h0);
  reg [(5'h17):(1'h0)] reg722 = (1'h0);
  reg [(5'h11):(1'h0)] reg723 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg725 = (1'h0);
  reg [(5'h18):(1'h0)] reg727 = (1'h0);
  reg [(5'h10):(1'h0)] reg730 = (1'h0);
  reg [(5'h17):(1'h0)] reg734 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg739 = (1'h0);
  reg [(5'h13):(1'h0)] reg740 = (1'h0);
  reg [(3'h4):(1'h0)] reg741 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg737 = (1'h0);
  reg [(5'h15):(1'h0)] reg743 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg746 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg747 = (1'h0);
  reg [(5'h16):(1'h0)] reg748 = (1'h0);
  reg [(5'h14):(1'h0)] reg749 = (1'h0);
  reg [(3'h7):(1'h0)] reg755 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg765 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg771 = (1'h0);
  reg [(5'h14):(1'h0)] reg772 = (1'h0);
  reg [(3'h4):(1'h0)] reg776 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg876 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg879 = (1'h0);
  reg [(5'h11):(1'h0)] reg880 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg883 = (1'h0);
  reg [(5'h11):(1'h0)] reg887 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg888 = (1'h0);
  reg [(5'h11):(1'h0)] reg891 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg892 = (1'h0);
  reg [(5'h12):(1'h0)] reg898 = (1'h0);
  reg [(4'he):(1'h0)] reg899 = (1'h0);
  reg [(5'h18):(1'h0)] reg902 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg904 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg905 = (1'h0);
  reg [(4'hd):(1'h0)] reg907 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg908 = (1'h0);
  reg [(4'hc):(1'h0)] reg914 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg918 = (1'h0);
  reg signed [(4'he):(1'h0)] reg919 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg920 = (1'h0);
  reg [(2'h2):(1'h0)] reg922 = (1'h0);
  reg [(3'h6):(1'h0)] reg923 = (1'h0);
  reg [(4'ha):(1'h0)] reg924 = (1'h0);
  reg [(3'h7):(1'h0)] reg930 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg931 = (1'h0);
  reg [(3'h5):(1'h0)] reg932 = (1'h0);
  reg [(4'ha):(1'h0)] reg933 = (1'h0);
  reg [(4'he):(1'h0)] reg935 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg936 = (1'h0);
  reg [(3'h4):(1'h0)] reg1140 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1141 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1425 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1423 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1420 = (1'h0);
  reg [(3'h7):(1'h0)] reg1419 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1414 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1411 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1410 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1409 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1406 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1404 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1403 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1400 = (1'h0);
  reg [(4'hf):(1'h0)] reg1399 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1396 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1395 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1382 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1391 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1389 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1387 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1385 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1384 = (1'h0);
  reg [(4'hc):(1'h0)] reg1383 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1382 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1379 = (1'h0);
  reg [(5'h16):(1'h0)] reg1378 = (1'h0);
  reg [(5'h18):(1'h0)] reg1377 = (1'h0);
  reg [(4'hf):(1'h0)] reg1375 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1372 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1369 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1367 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1366 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1360 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1359 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1357 = (1'h0);
  reg [(4'h8):(1'h0)] reg1356 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1354 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1352 = (1'h0);
  reg [(4'hd):(1'h0)] reg1348 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1347 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1346 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1344 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1343 = (1'h0);
  reg [(4'he):(1'h0)] reg1342 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1341 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1340 = (1'h0);
  reg [(3'h7):(1'h0)] reg1339 = (1'h0);
  reg [(5'h16):(1'h0)] reg934 = (1'h0);
  reg [(3'h5):(1'h0)] forvar927 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg926 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg929 = (1'h0);
  reg [(5'h14):(1'h0)] reg928 = (1'h0);
  reg [(3'h4):(1'h0)] reg927 = (1'h0);
  reg [(4'h9):(1'h0)] forvar926 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg925 = (1'h0);
  reg [(4'hc):(1'h0)] forvar921 = (1'h0);
  reg [(4'h8):(1'h0)] forvar917 = (1'h0);
  reg [(5'h18):(1'h0)] forvar916 = (1'h0);
  reg [(2'h3):(1'h0)] forvar905 = (1'h0);
  reg [(2'h3):(1'h0)] reg915 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg913 = (1'h0);
  reg [(5'h17):(1'h0)] reg912 = (1'h0);
  reg [(4'h9):(1'h0)] reg911 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar910 = (1'h0);
  reg [(4'h9):(1'h0)] reg909 = (1'h0);
  reg [(3'h7):(1'h0)] reg906 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg901 = (1'h0);
  reg [(4'hf):(1'h0)] forvar900 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar895 = (1'h0);
  reg [(3'h5):(1'h0)] reg897 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg896 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg895 = (1'h0);
  reg [(4'hb):(1'h0)] reg894 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg893 = (1'h0);
  reg [(5'h17):(1'h0)] reg890 = (1'h0);
  reg [(5'h14):(1'h0)] forvar889 = (1'h0);
  reg [(4'hb):(1'h0)] reg886 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar885 = (1'h0);
  reg [(3'h7):(1'h0)] forvar877 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg884 = (1'h0);
  reg [(5'h15):(1'h0)] reg882 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg881 = (1'h0);
  reg [(4'ha):(1'h0)] reg878 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg877 = (1'h0);
  reg [(5'h11):(1'h0)] reg875 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg874 = (1'h0);
  reg [(5'h15):(1'h0)] reg777 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar775 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg774 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg773 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg770 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg769 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar768 = (1'h0);
  reg [(5'h17):(1'h0)] reg767 = (1'h0);
  reg [(4'hd):(1'h0)] forvar766 = (1'h0);
  reg [(5'h12):(1'h0)] reg764 = (1'h0);
  reg [(4'hf):(1'h0)] reg763 = (1'h0);
  reg [(4'ha):(1'h0)] reg762 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg761 = (1'h0);
  reg [(5'h12):(1'h0)] reg760 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar759 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg758 = (1'h0);
  reg [(4'hc):(1'h0)] reg757 = (1'h0);
  reg [(5'h11):(1'h0)] reg756 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg754 = (1'h0);
  reg [(3'h4):(1'h0)] reg753 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar752 = (1'h0);
  reg [(5'h13):(1'h0)] reg751 = (1'h0);
  reg [(5'h11):(1'h0)] reg750 = (1'h0);
  reg [(5'h11):(1'h0)] reg745 = (1'h0);
  reg [(2'h3):(1'h0)] forvar744 = (1'h0);
  reg [(3'h7):(1'h0)] reg742 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar734 = (1'h0);
  reg [(3'h6):(1'h0)] reg738 = (1'h0);
  reg [(4'he):(1'h0)] forvar737 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg736 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg735 = (1'h0);
  reg [(4'he):(1'h0)] reg733 = (1'h0);
  reg [(5'h14):(1'h0)] reg732 = (1'h0);
  reg [(4'hf):(1'h0)] reg731 = (1'h0);
  reg [(4'he):(1'h0)] reg729 = (1'h0);
  reg [(5'h10):(1'h0)] reg728 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg726 = (1'h0);
  reg [(5'h13):(1'h0)] forvar722 = (1'h0);
  reg [(4'hd):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg720 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg719 = (1'h0);
  reg [(3'h6):(1'h0)] reg717 = (1'h0);
  reg [(3'h4):(1'h0)] reg716 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg714 = (1'h0);
  reg [(4'h8):(1'h0)] reg713 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg711 = (1'h0);
  reg [(5'h13):(1'h0)] reg710 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar701 = (1'h0);
  reg [(4'hf):(1'h0)] reg709 = (1'h0);
  reg [(4'hb):(1'h0)] forvar707 = (1'h0);
  reg [(4'hc):(1'h0)] reg706 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg705 = (1'h0);
  reg signed [(4'he):(1'h0)] reg700 = (1'h0);
  reg [(4'hb):(1'h0)] reg699 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg698 = (1'h0);
  reg [(4'he):(1'h0)] reg695 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg692 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg690 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg689 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg687 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg685 = (1'h0);
  assign y = {wire1595,
                 wire1593,
                 wire1431,
                 wire1337,
                 wire1335,
                 wire1138,
                 wire872,
                 reg1596,
                 reg1430,
                 reg1429,
                 reg1428,
                 reg1427,
                 reg1426,
                 reg1424,
                 reg1422,
                 reg1421,
                 reg1414,
                 reg1418,
                 reg1417,
                 reg1416,
                 reg1415,
                 reg1413,
                 reg1400,
                 reg1396,
                 reg1412,
                 reg1408,
                 reg1407,
                 reg1405,
                 reg1402,
                 reg1401,
                 reg1398,
                 reg1397,
                 reg1394,
                 reg1393,
                 reg1392,
                 reg1390,
                 reg1388,
                 reg1386,
                 reg1381,
                 reg1380,
                 reg1376,
                 reg1374,
                 reg1373,
                 reg1371,
                 reg1370,
                 reg1368,
                 reg1365,
                 reg1364,
                 reg1363,
                 reg1362,
                 reg1361,
                 reg1358,
                 reg1355,
                 reg1353,
                 reg1351,
                 reg1350,
                 reg1349,
                 reg1345,
                 reg1338,
                 reg686,
                 reg688,
                 reg691,
                 reg693,
                 reg694,
                 reg696,
                 reg697,
                 reg701,
                 reg702,
                 reg703,
                 reg704,
                 reg708,
                 reg707,
                 reg712,
                 reg715,
                 reg718,
                 reg721,
                 reg722,
                 reg723,
                 reg725,
                 reg727,
                 reg730,
                 reg734,
                 reg739,
                 reg740,
                 reg741,
                 reg737,
                 reg743,
                 reg746,
                 reg747,
                 reg748,
                 reg749,
                 reg755,
                 reg765,
                 reg771,
                 reg772,
                 reg776,
                 reg876,
                 reg879,
                 reg880,
                 reg883,
                 reg887,
                 reg888,
                 reg891,
                 reg892,
                 reg898,
                 reg899,
                 reg902,
                 reg904,
                 reg905,
                 reg907,
                 reg908,
                 reg914,
                 reg918,
                 reg919,
                 reg920,
                 reg922,
                 reg923,
                 reg924,
                 reg930,
                 reg931,
                 reg932,
                 reg933,
                 reg935,
                 reg936,
                 reg1140,
                 reg1141,
                 forvar1425,
                 reg1423,
                 forvar1420,
                 reg1419,
                 forvar1414,
                 reg1411,
                 reg1410,
                 forvar1409,
                 reg1406,
                 reg1404,
                 reg1403,
                 forvar1400,
                 reg1399,
                 forvar1396,
                 reg1395,
                 reg1382,
                 forvar1391,
                 reg1389,
                 reg1387,
                 forvar1385,
                 reg1384,
                 reg1383,
                 forvar1382,
                 forvar1379,
                 reg1378,
                 reg1377,
                 reg1375,
                 forvar1372,
                 forvar1369,
                 reg1367,
                 forvar1366,
                 forvar1360,
                 forvar1359,
                 forvar1357,
                 reg1356,
                 reg1354,
                 forvar1352,
                 reg1348,
                 reg1347,
                 reg1346,
                 reg1344,
                 reg1343,
                 reg1342,
                 forvar1341,
                 forvar1340,
                 reg1339,
                 reg934,
                 forvar927,
                 reg926,
                 reg929,
                 reg928,
                 reg927,
                 forvar926,
                 reg925,
                 forvar921,
                 forvar917,
                 forvar916,
                 forvar905,
                 reg915,
                 reg913,
                 reg912,
                 reg911,
                 forvar910,
                 reg909,
                 reg906,
                 reg903,
                 reg901,
                 forvar900,
                 forvar895,
                 reg897,
                 reg896,
                 reg895,
                 reg894,
                 reg893,
                 reg890,
                 forvar889,
                 reg886,
                 forvar885,
                 forvar877,
                 reg884,
                 reg882,
                 reg881,
                 reg878,
                 reg877,
                 reg875,
                 reg874,
                 reg777,
                 forvar775,
                 reg774,
                 reg773,
                 reg770,
                 reg769,
                 forvar768,
                 reg767,
                 forvar766,
                 reg764,
                 reg763,
                 reg762,
                 reg761,
                 reg760,
                 forvar759,
                 reg758,
                 reg757,
                 reg756,
                 reg754,
                 reg753,
                 forvar752,
                 reg751,
                 reg750,
                 reg745,
                 forvar744,
                 reg742,
                 forvar734,
                 reg738,
                 forvar737,
                 reg736,
                 reg735,
                 reg733,
                 reg732,
                 reg731,
                 reg729,
                 reg728,
                 reg726,
                 forvar722,
                 reg724,
                 reg720,
                 reg719,
                 reg717,
                 reg716,
                 reg714,
                 reg713,
                 reg711,
                 reg710,
                 forvar701,
                 reg709,
                 forvar707,
                 reg706,
                 reg705,
                 reg700,
                 reg699,
                 reg698,
                 reg695,
                 reg692,
                 reg690,
                 reg689,
                 reg687,
                 reg685,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg685 = ($unsigned((-((wire682 ?
          wire680 : wire680) - wire680[(3'h7):(1'h1)]))) + (8'ha3));
      if (({{(8'h9d), wire680}, (wire681 < $unsigned($unsigned(wire683)))} ?
          wire684[(5'h11):(4'hf)] : wire680))
        begin
          reg686 <= ($unsigned((+wire683)) ?
              wire683[(4'hb):(4'hb)] : (($unsigned($signed(wire682)) != $signed((wire682 ?
                  wire683 : wire684))) != (!((wire680 ?
                  wire680 : wire682) <<< wire680))));
          if (((8'ha8) ?
              (wire684[(3'h5):(2'h2)] ?
                  $signed((~&((7'h42) > wire683))) : {wire683}) : (wire681 > wire680)))
            begin
              reg687 = (|({{$signed(wire682), (|wire680)},
                  $unsigned($unsigned(reg685))} > $unsigned(((^~wire681) <<< $unsigned(wire684)))));
              reg688 <= $signed((-$unsigned(reg685[(3'h4):(1'h1)])));
              reg689 = wire683;
              reg690 = (-($signed(((reg686 || reg689) ?
                  {reg689, reg687} : $unsigned(wire680))) == reg685));
              reg691 <= $signed((~^{reg685[(1'h1):(1'h1)]}));
            end
          else
            begin
              reg687 = $unsigned(wire682);
              reg689 = $unsigned($signed((reg686 ^~ ((|reg687) ?
                  ((8'hbc) != (8'ha6)) : $unsigned(wire680)))));
              reg690 = ((~(!((+wire681) | $signed(reg686)))) ?
                  ($signed(((wire682 ?
                      wire684 : wire684) || $signed(reg690))) | reg687[(2'h2):(2'h2)]) : wire680);
            end
          reg692 = (~&reg688);
          if ($unsigned(reg685[(3'h6):(3'h6)]))
            begin
              reg693 <= wire680[(3'h5):(3'h4)];
              reg694 <= ((((wire683 ? (~|reg685) : reg693) ?
                      ((^reg687) ?
                          (wire683 << reg688) : $signed(wire682)) : (^(reg691 * (8'haa)))) << reg686) ?
                  (7'h40) : reg688[(1'h0):(1'h0)]);
              reg695 = $unsigned(($signed(reg691) ?
                  reg691[(5'h12):(2'h3)] : reg690[(1'h0):(1'h0)]));
              reg696 <= reg688;
              reg697 <= (($unsigned(reg685) ?
                  $signed($signed(wire680[(4'h9):(1'h0)])) : {reg686[(3'h4):(1'h0)]}) >>> $signed(((reg695 || reg688) ?
                  (&$signed(reg686)) : ({wire684} < reg693))));
            end
          else
            begin
              reg693 <= reg686[(2'h3):(2'h2)];
              reg694 <= ({$unsigned(({reg696, reg688} & $unsigned(wire684)))} ?
                  reg686[(2'h2):(1'h1)] : $unsigned(reg696));
              reg696 <= reg697[(3'h7):(1'h1)];
              reg698 = ((((&(~&reg690)) >= (^(|(8'h9e)))) ?
                      reg689 : (&$unsigned(wire681))) ?
                  (+{{((8'hba) >= reg687), ((7'h4a) ? reg685 : wire681)},
                      ((reg697 ?
                          reg696 : (7'h42)) * $unsigned((8'hb0)))}) : (reg685[(1'h0):(1'h0)] >>> (($unsigned(reg688) * $signed(reg685)) ?
                      $signed(reg695[(1'h0):(1'h0)]) : reg696)));
              reg699 = $signed((~(reg695 ? {(-reg697)} : $unsigned(reg689))));
            end
          reg700 = wire680;
        end
      else
        begin
          reg687 = (8'hbf);
        end
    end
  always
    @(posedge clk) begin
      if (wire684[(5'h13):(1'h0)])
        begin
          reg701 <= ((-wire683[(2'h2):(2'h2)]) ?
              (!((8'h9f) ?
                  reg686[(3'h4):(1'h1)] : (reg693[(1'h1):(1'h0)] ^~ ((7'h4a) ?
                      reg694 : reg696)))) : ($signed(((&reg697) >> (reg686 + reg686))) ?
                  (!{wire680,
                      wire683[(3'h4):(1'h0)]}) : $unsigned(($signed(wire684) ^ (wire682 ?
                      wire684 : reg694)))));
          if ((reg697[(1'h1):(1'h0)] * ((~$unsigned((wire684 ?
              reg686 : reg691))) == $signed((!(reg691 ? wire684 : reg693))))))
            begin
              reg702 <= reg701;
              reg703 <= reg686;
              reg704 <= (~^$unsigned(($signed((reg696 < reg696)) ?
                  reg697[(4'h9):(4'h9)] : reg703[(3'h5):(2'h3)])));
              reg705 = $unsigned($unsigned((reg704[(2'h3):(1'h1)] ?
                  ((8'ha8) < (reg694 != (8'hb2))) : {$signed(reg694)})));
            end
          else
            begin
              reg702 <= $unsigned((+$unsigned(reg688)));
              reg703 <= $unsigned((reg704 == (~^(8'h9f))));
              reg704 <= reg693;
            end
          reg706 = $signed((&wire682));
          for (forvar707 = (1'h0); (forvar707 < (1'h1)); forvar707 = (forvar707 + (1'h1)))
            begin
              reg708 <= reg702;
            end
          reg709 = ((reg701[(4'hc):(3'h5)] ?
              $signed(reg705) : $unsigned(reg686[(1'h0):(1'h0)])) ^ reg688);
        end
      else
        begin
          for (forvar701 = (1'h0); (forvar701 < (3'h4)); forvar701 = (forvar701 + (1'h1)))
            begin
              reg705 = reg708;
              reg707 <= $unsigned(wire683);
              reg709 = reg707[(1'h1):(1'h1)];
            end
          reg710 = {reg703};
          if ($signed(reg701))
            begin
              reg711 = {(8'hb7), reg686[(3'h4):(2'h3)]};
              reg712 <= (reg688[(4'hb):(2'h2)] < ((({wire681} <<< $signed(reg710)) | $unsigned(reg711)) || {(forvar701 | reg693),
                  ((reg703 ? reg704 : wire683) ^~ $signed(reg701))}));
              reg713 = (~^(~{reg686[(1'h1):(1'h0)]}));
            end
          else
            begin
              reg711 = (|(!((+$signed(reg686)) >= (reg707[(1'h0):(1'h0)] != $signed(reg694)))));
            end
          if (reg688)
            begin
              reg714 = (~&{($unsigned($unsigned(reg686)) >= reg712),
                  reg712[(3'h4):(2'h3)]});
              reg715 <= forvar707[(4'ha):(2'h2)];
              reg716 = (wire680 ^ reg714[(1'h1):(1'h0)]);
              reg717 = (&((((wire684 ? wire680 : reg688) ?
                  reg713[(2'h2):(2'h2)] : {reg701,
                      forvar701}) && reg706) < wire681[(4'ha):(2'h2)]));
            end
          else
            begin
              reg714 = (&((^(8'haf)) ? reg713 : reg704));
              reg716 = reg707;
              reg718 <= reg703;
            end
        end
      if ((~$signed(((~^(reg694 ? wire682 : reg705)) ?
          $signed(reg709[(3'h7):(3'h4)]) : (&$unsigned(reg706))))))
        begin
          if ((((reg711 ?
              $signed((reg696 ?
                  forvar701 : reg697)) : $unsigned((~|reg713))) + $signed(wire682)) <<< (($signed($signed(reg716)) ^~ {$unsigned((8'h9d)),
                  (reg713 ? reg701 : reg707)}) ?
              reg714[(2'h3):(2'h2)] : $signed({$signed(reg705)}))))
            begin
              reg719 = reg691;
              reg720 = (reg708 & $signed(reg694[(3'h4):(1'h1)]));
              reg721 <= $unsigned(reg694[(1'h0):(1'h0)]);
              reg722 <= ($unsigned(wire681[(3'h5):(2'h3)]) * reg711);
              reg723 <= reg706[(3'h5):(2'h2)];
            end
          else
            begin
              reg719 = (|((reg706 ?
                      reg694[(3'h7):(3'h4)] : $unsigned(reg721[(4'he):(4'h8)])) ?
                  (&$unsigned(((8'haa) ? reg709 : wire680))) : (reg708 ?
                      {$unsigned(wire681),
                          (reg704 ? reg715 : wire682)} : $unsigned((reg722 ?
                          reg713 : wire684)))));
              reg721 <= $unsigned({wire680[(1'h1):(1'h0)]});
              reg722 <= (~^(reg715 ?
                  (&reg696[(2'h2):(1'h0)]) : (|($unsigned(reg688) && reg722))));
              reg724 = reg688[(4'he):(2'h2)];
            end
        end
      else
        begin
          reg721 <= $signed((~&($signed((reg724 ? reg724 : reg716)) ?
              $unsigned(wire681) : reg688)));
          for (forvar722 = (1'h0); (forvar722 < (2'h3)); forvar722 = (forvar722 + (1'h1)))
            begin
              reg723 <= {$signed(($signed($signed(reg710)) | $signed((!reg708))))};
            end
          reg725 <= $unsigned(reg715);
          reg726 = $unsigned(reg711);
          if (($signed((-((forvar701 >= reg702) ?
                  $signed(reg714) : (reg717 ^ reg686)))) ?
              reg717 : ($signed((8'h9d)) - (reg704[(4'hc):(3'h7)] ?
                  {{reg724}, $unsigned(reg707)} : {forvar701[(3'h6):(3'h4)],
                      (reg706 ^ (8'ha7))}))))
            begin
              reg727 <= ($unsigned((~($unsigned((8'ha1)) & $unsigned(reg707)))) || reg714);
              reg728 = $signed($signed(reg712));
              reg729 = $unsigned($signed((reg724[(3'h5):(3'h4)] ?
                  ((reg714 >>> forvar707) >= $signed(reg697)) : reg727)));
            end
          else
            begin
              reg727 <= $unsigned((reg725 ?
                  reg723[(4'hd):(3'h6)] : (reg721 >>> {(reg724 - reg703)})));
              reg728 = $unsigned(reg703);
              reg730 <= (|(forvar701[(2'h3):(1'h1)] ? reg721 : reg686));
              reg731 = (|reg694[(4'hb):(3'h4)]);
              reg732 = ($signed((~|{(&reg731),
                  $signed(forvar722)})) <<< reg703);
            end
        end
      reg733 = ((($signed($signed(reg732)) << {wire680[(1'h1):(1'h1)],
          $signed(reg727)}) > {(-reg721[(4'h9):(2'h2)]),
          (~^reg703)}) ~^ reg729[(4'h9):(4'h8)]);
      if (((8'ha9) ?
          ((7'h40) ?
              (($signed(reg704) ? (reg720 <= wire684) : $signed(forvar722)) ?
                  reg726[(1'h0):(1'h0)] : ((reg693 >= (8'had)) ?
                      (reg723 ?
                          reg693 : reg713) : (wire682 << reg710))) : (reg686[(2'h3):(2'h2)] != forvar707[(3'h7):(3'h4)])) : ((reg709[(4'hd):(4'h8)] >= (((7'h43) ?
              wire683 : reg703) & wire683[(5'h12):(4'ha)])) >>> reg703[(1'h1):(1'h1)])))
        begin
          reg734 <= reg716;
          reg735 = (8'hac);
          reg736 = ($unsigned({reg694}) <<< reg723[(3'h5):(3'h4)]);
          for (forvar737 = (1'h0); (forvar737 < (2'h2)); forvar737 = (forvar737 + (1'h1)))
            begin
              reg738 = ($unsigned($unsigned($signed($unsigned(reg736)))) ~^ (|wire684[(4'hd):(3'h6)]));
              reg739 <= $signed((!forvar722[(1'h0):(1'h0)]));
              reg740 <= $signed($signed(reg735[(3'h5):(1'h1)]));
              reg741 <= $signed($signed((reg693 ?
                  reg733 : (~^(reg708 ? reg718 : reg731)))));
            end
        end
      else
        begin
          for (forvar734 = (1'h0); (forvar734 < (2'h2)); forvar734 = (forvar734 + (1'h1)))
            begin
              reg737 <= {((reg741[(1'h0):(1'h0)] ?
                          $signed((&reg703)) : $signed((|(8'ha3)))) ?
                      reg696 : {{((8'hb3) - forvar737), (reg711 >>> reg734)}}),
                  (^$unsigned(reg703[(1'h0):(1'h0)]))};
              reg739 <= ((~reg707[(1'h1):(1'h1)]) >>> $signed(reg741[(2'h3):(2'h2)]));
              reg740 <= ((-reg735) ? (!reg719) : reg712[(4'h8):(3'h7)]);
              reg742 = (reg713[(4'h8):(1'h0)] * reg714[(1'h0):(1'h0)]);
            end
          reg743 <= $signed($signed($signed(((reg733 ?
              (8'hae) : reg686) & {(7'h46)}))));
          for (forvar744 = (1'h0); (forvar744 < (3'h4)); forvar744 = (forvar744 + (1'h1)))
            begin
              reg745 = reg725[(1'h0):(1'h0)];
            end
          reg746 <= reg717[(1'h0):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      reg747 <= wire681[(3'h7):(1'h1)];
      reg748 <= reg718;
      reg749 <= reg746[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg750 = $signed(((8'ha9) ? reg686[(2'h3):(2'h3)] : $signed(reg727)));
      reg751 = $signed(reg704);
      for (forvar752 = (1'h0); (forvar752 < (2'h3)); forvar752 = (forvar752 + (1'h1)))
        begin
          reg753 = ((8'hbc) ?
              $signed($signed(reg727[(4'hf):(3'h4)])) : ((8'h9e) ?
                  $unsigned(wire681[(1'h1):(1'h0)]) : ($signed({(8'hb0)}) ?
                      reg686 : reg702)));
          if ($signed(reg691[(3'h5):(1'h1)]))
            begin
              reg754 = $signed((((reg694 ? (reg747 * reg753) : (!reg750)) ?
                      ($signed(wire681) <<< $unsigned(wire684)) : {(^~wire681),
                          {wire682, reg715}}) ?
                  reg697 : reg708));
              reg755 <= reg741[(1'h1):(1'h1)];
              reg756 = $unsigned(reg715[(1'h0):(1'h0)]);
              reg757 = $signed((({$signed(reg739), $signed(reg750)} ?
                  ($unsigned((8'ha5)) ?
                      (^wire680) : $unsigned((8'ha7))) : (~|$unsigned(reg702))) <<< reg737[(4'hf):(4'hd)]));
              reg758 = (&$signed((~|$unsigned(forvar752))));
            end
          else
            begin
              reg754 = $unsigned($unsigned(reg725));
            end
          for (forvar759 = (1'h0); (forvar759 < (1'h0)); forvar759 = (forvar759 + (1'h1)))
            begin
              reg760 = reg707;
              reg761 = {(((~^forvar752[(5'h12):(2'h2)]) & ((reg707 ?
                          reg758 : reg708) ?
                      ((8'h9f) & reg757) : reg750)) ^ ($signed((reg697 >> reg722)) ?
                      (~^wire681[(4'ha):(4'ha)]) : reg691[(1'h1):(1'h0)]))};
              reg762 = (wire681[(2'h3):(2'h3)] + {$signed(reg722[(1'h0):(1'h0)])});
              reg763 = ($unsigned({(-$signed(reg715)),
                  $signed($signed(reg750))}) >> (!reg746));
              reg764 = $signed((~|reg753[(2'h2):(2'h2)]));
            end
        end
      reg765 <= ((8'hbd) - (^reg746));
      for (forvar766 = (1'h0); (forvar766 < (1'h0)); forvar766 = (forvar766 + (1'h1)))
        begin
          reg767 = reg696[(1'h0):(1'h0)];
          for (forvar768 = (1'h0); (forvar768 < (3'h4)); forvar768 = (forvar768 + (1'h1)))
            begin
              reg769 = {{$signed(reg694[(1'h1):(1'h1)])}};
              reg770 = ($unsigned((|$signed($unsigned(forvar768)))) ?
                  ({(!$signed(wire682)), reg688} ?
                      reg693 : {forvar759[(4'hc):(1'h0)],
                          (reg701[(2'h2):(1'h0)] ?
                              reg730[(4'h9):(3'h4)] : $unsigned(reg747))}) : {reg753});
              reg771 <= ((((^reg737) <= (^(~^reg762))) <<< ($unsigned(reg727[(5'h16):(5'h14)]) << (|(reg756 ?
                  reg697 : reg691)))) <<< (8'hbc));
              reg772 <= $signed($unsigned(forvar759[(1'h1):(1'h1)]));
              reg773 = $unsigned((reg769 ?
                  (((reg693 >> reg712) ?
                          $unsigned(wire680) : reg740[(4'h8):(1'h1)]) ?
                      ($signed(reg734) | (reg703 - reg697)) : ((reg741 ?
                          (8'h9f) : reg767) & (reg767 << reg748))) : ((reg763 ?
                          $unsigned((8'hb7)) : reg772) ?
                      $unsigned((!(8'hb8))) : reg749[(4'h8):(4'h8)])));
            end
          reg774 = $signed($unsigned($unsigned($unsigned($signed(reg727)))));
          for (forvar775 = (1'h0); (forvar775 < (2'h3)); forvar775 = (forvar775 + (1'h1)))
            begin
              reg776 <= (((((reg727 ? wire681 : reg722) ^~ ((8'hae) ?
                          reg725 : wire681)) >> reg773[(3'h6):(3'h5)]) ?
                      reg737 : reg722[(4'ha):(4'h9)]) ?
                  (((^$unsigned(wire682)) >> $unsigned((reg743 ?
                      reg751 : reg723))) != {{$signed(reg737)},
                      ((^~reg749) ~^ {(8'ha4), reg704})}) : $signed((8'ha9)));
              reg777 = (8'hbb);
            end
        end
    end
  module778 #() modinst873 (wire872, clk, reg703, reg734, reg740, wire684, reg746);
  always
    @(posedge clk) begin
      reg874 = {{$unsigned(reg734),
              $unsigned(((reg721 ? reg697 : reg741) ?
                  (&reg703) : reg740[(4'he):(4'he)]))}};
      if (reg730)
        begin
          reg875 = reg755[(3'h5):(2'h3)];
          reg876 <= (|(($signed(reg704) ^ ((reg776 ?
                  reg755 : reg772) >= (reg715 ^~ reg765))) ?
              {$signed((reg739 != reg748)),
                  ((reg874 ? reg723 : reg718) || {reg772,
                      reg718})} : (wire684 ^ reg697[(2'h3):(2'h2)])));
          if ((~^($unsigned((reg722 ? reg715 : $signed(reg702))) ?
              (reg686 ? wire872 : $unsigned(reg704)) : reg712[(4'hf):(4'ha)])))
            begin
              reg877 = $signed((((reg688 + (reg776 & wire681)) ?
                      reg701[(2'h3):(2'h2)] : reg748[(4'he):(1'h0)]) ?
                  (-reg704[(4'hc):(2'h3)]) : $signed($signed($signed(reg737)))));
              reg878 = reg691;
            end
          else
            begin
              reg879 <= (((reg776 ?
                      ({reg701, (8'ha9)} == (^reg877)) : ((reg722 ?
                          reg737 : reg741) | reg693[(3'h4):(2'h2)])) + (((reg737 && wire680) ?
                          (+reg712) : reg765) ?
                      reg748[(2'h2):(1'h1)] : (8'hae))) ?
                  ($unsigned($signed(reg749)) ?
                      $signed((~&reg688[(5'h14):(4'ha)])) : ($unsigned(reg723[(3'h5):(1'h1)]) ?
                          $signed((reg875 ?
                              reg703 : reg737)) : reg876)) : $unsigned((+($signed(reg776) > $unsigned(reg704)))));
              reg880 <= ($signed((reg701[(4'hc):(1'h0)] ~^ (reg765[(4'hd):(1'h0)] ?
                  reg715 : ((8'ha2) > (7'h45))))) - (reg691[(1'h1):(1'h1)] ?
                  (reg725[(2'h2):(2'h2)] >> $unsigned(reg875)) : ($signed(reg765[(4'h8):(3'h7)]) ?
                      $signed(reg772) : {{reg694}})));
              reg881 = ($unsigned((~&$signed((reg701 | wire681)))) - ($unsigned(($unsigned((8'h9e)) ?
                      {reg704, reg697} : reg743)) ?
                  {((reg691 ?
                          (7'h42) : reg702) << reg749)} : ((~&$signed(reg879)) - {$signed((8'ha0))})));
              reg882 = ((({$unsigned(wire682), {reg727}} ?
                          (-reg730[(4'he):(4'ha)]) : {reg718[(4'h9):(4'h8)]}) ?
                      $unsigned((reg715 ?
                          reg727[(1'h0):(1'h0)] : $unsigned(reg881))) : {reg712[(2'h3):(2'h2)]}) ?
                  (($unsigned($signed(wire680)) <<< reg703) <<< (($unsigned(reg721) <<< ((8'h9c) ?
                          reg741 : reg740)) ?
                      $signed({reg702}) : $signed((reg703 ?
                          wire681 : reg715)))) : $signed(reg876));
            end
          reg883 <= $signed((&(+(8'hb0))));
          reg884 = reg776[(3'h4):(2'h2)];
        end
      else
        begin
          reg876 <= {wire681[(4'h8):(3'h4)]};
          for (forvar877 = (1'h0); (forvar877 < (2'h2)); forvar877 = (forvar877 + (1'h1)))
            begin
              reg879 <= (reg737[(4'hf):(4'h9)] ?
                  reg725[(1'h1):(1'h0)] : wire681[(1'h1):(1'h0)]);
              reg880 <= $unsigned($signed((((reg739 ? reg741 : reg701) ?
                  reg883[(3'h4):(3'h4)] : $signed(reg707)) * (+$signed(reg712)))));
            end
          if ((($unsigned((8'hbe)) ?
              $signed(reg772[(4'h8):(2'h3)]) : ({(^reg707), reg772} ?
                  reg686 : (((7'h43) >>> forvar877) || $unsigned(reg737)))) & {(($unsigned(reg877) ?
                      {reg707, (8'ha4)} : ((8'ha0) && reg696)) ?
                  reg688[(4'h8):(3'h4)] : ({(8'had), (8'hbd)} ?
                      reg686 : {reg725})),
              reg688}))
            begin
              reg883 <= ($unsigned((($unsigned(reg765) && (8'hbd)) * {$unsigned((8'hb9)),
                  (reg688 | reg879)})) - reg712);
            end
          else
            begin
              reg881 = $unsigned($unsigned($unsigned(($unsigned(reg701) << {reg740,
                  reg776}))));
              reg882 = (reg730 ?
                  (reg697 ?
                      ($unsigned((~&reg693)) || ($signed(reg701) ?
                          $signed(reg701) : ((7'h47) ?
                              wire680 : reg884))) : (({reg881,
                          reg704} << (reg882 ?
                          reg723 : reg743)) << reg746[(2'h2):(2'h2)])) : ((^reg776) >> (wire684 ?
                      reg874[(4'h9):(3'h6)] : (reg688[(4'hd):(1'h0)] ~^ $signed(reg771)))));
              reg884 = reg722;
            end
        end
      for (forvar885 = (1'h0); (forvar885 < (2'h2)); forvar885 = (forvar885 + (1'h1)))
        begin
          reg886 = reg875[(4'h8):(3'h5)];
          reg887 <= (~(~&$signed((7'h45))));
          reg888 <= $signed(((reg765[(2'h3):(2'h2)] ?
                  $signed((8'hb7)) : reg721[(4'hf):(4'he)]) ?
              ($unsigned($unsigned(reg881)) ?
                  {reg876} : reg727[(4'hf):(4'hd)]) : (((reg702 ?
                      reg739 : reg707) ?
                  {reg696} : (reg702 ?
                      reg743 : reg877)) ^ reg886[(2'h3):(2'h3)])));
          for (forvar889 = (1'h0); (forvar889 < (3'h4)); forvar889 = (forvar889 + (1'h1)))
            begin
              reg890 = ((7'h47) ?
                  {{($signed((8'h9f)) >>> reg694[(1'h0):(1'h0)])}} : wire681);
              reg891 <= reg725;
              reg892 <= reg771;
              reg893 = ((&reg730[(3'h4):(1'h0)]) || reg694);
            end
        end
      reg894 = reg701[(4'hf):(4'h8)];
      if ((reg892 < $unsigned($signed(reg691))))
        begin
          if ((+((~&((reg772 >>> reg746) ? (|reg748) : {reg730})) ?
              (((&reg893) >> $signed(reg694)) ?
                  reg701 : $unsigned($unsigned(reg743))) : $signed(reg894[(4'h8):(3'h7)]))))
            begin
              reg895 = (+reg892);
              reg896 = (((reg739[(1'h0):(1'h0)] == {reg688,
                      reg703[(2'h2):(1'h0)]}) ?
                  ($signed((&reg893)) - (((7'h45) ?
                      (7'h44) : reg715) <<< reg765[(3'h6):(3'h6)])) : wire684) < $unsigned({{$unsigned(reg697)},
                  ((^~forvar885) ? (~^wire684) : $signed(forvar877))}));
              reg897 = $unsigned(($signed(reg892[(2'h3):(1'h1)]) + (reg701 ^~ reg755[(1'h1):(1'h1)])));
            end
          else
            begin
              reg895 = reg725[(2'h3):(2'h2)];
            end
        end
      else
        begin
          for (forvar895 = (1'h0); (forvar895 < (1'h1)); forvar895 = (forvar895 + (1'h1)))
            begin
              reg898 <= $unsigned((!($unsigned($unsigned(reg723)) ?
                  (~|(8'hb0)) : $unsigned((reg743 ? reg740 : (8'hae))))));
            end
          reg899 <= $unsigned((&reg897[(3'h5):(1'h0)]));
          for (forvar900 = (1'h0); (forvar900 < (2'h2)); forvar900 = (forvar900 + (1'h1)))
            begin
              reg901 = reg776;
              reg902 <= ($signed((reg884[(2'h2):(1'h0)] <<< $unsigned(wire684))) >= reg896);
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed(reg746))
        begin
          if (reg715)
            begin
              reg903 = {reg730[(4'hb):(4'ha)]};
              reg904 <= (((($signed(reg776) ? {reg703} : (reg712 >= reg704)) ?
                      ((!reg883) != $unsigned(reg743)) : $signed($signed(reg887))) ?
                  (^$signed(reg696)) : $signed($unsigned(((8'hb9) ~^ reg898)))) & {reg693,
                  $unsigned(reg755)});
              reg905 <= (+(~({reg741} ?
                  reg883[(4'h8):(3'h7)] : ((wire684 >= reg718) ?
                      (reg904 > reg765) : (reg776 ? reg686 : wire872)))));
            end
          else
            begin
              reg903 = (~^($signed(reg725) && reg741));
              reg904 <= (^$unsigned((8'had)));
              reg906 = $unsigned(reg904[(1'h0):(1'h0)]);
              reg907 <= {($signed(reg715) > (($signed(reg888) < (reg892 ?
                          reg743 : (8'h9f))) ?
                      $unsigned($signed(reg734)) : $unsigned(reg718[(3'h4):(2'h2)]))),
                  (($unsigned({reg741}) ^ $signed(reg691[(5'h12):(2'h2)])) ?
                      reg755[(1'h0):(1'h0)] : reg708)};
              reg908 <= reg704[(4'hf):(4'hb)];
            end
          reg909 = $signed($signed(reg686[(3'h4):(1'h0)]));
          for (forvar910 = (1'h0); (forvar910 < (1'h0)); forvar910 = (forvar910 + (1'h1)))
            begin
              reg911 = (reg909[(3'h7):(2'h3)] < (reg727 ?
                  wire683 : reg739[(3'h4):(2'h3)]));
              reg912 = reg765;
              reg913 = $signed($signed(reg902));
              reg914 <= reg686;
            end
          reg915 = (8'h9e);
        end
      else
        begin
          reg904 <= reg701[(5'h12):(3'h5)];
          for (forvar905 = (1'h0); (forvar905 < (1'h1)); forvar905 = (forvar905 + (1'h1)))
            begin
              reg907 <= reg879;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar916 = (1'h0); (forvar916 < (1'h1)); forvar916 = (forvar916 + (1'h1)))
        begin
          for (forvar917 = (1'h0); (forvar917 < (1'h1)); forvar917 = (forvar917 + (1'h1)))
            begin
              reg918 <= $unsigned((^~({reg765[(5'h13):(4'hd)],
                      (reg691 >>> forvar916)} ?
                  reg740 : {(8'ha1), (8'hb0)})));
              reg919 <= $signed(reg771);
              reg920 <= $unsigned(reg686);
            end
          for (forvar921 = (1'h0); (forvar921 < (3'h4)); forvar921 = (forvar921 + (1'h1)))
            begin
              reg922 <= (reg727[(3'h7):(3'h7)] ?
                  (~^(&wire872[(1'h0):(1'h0)])) : (reg708 ^~ {(7'h47)}));
              reg923 <= (((^~reg686[(2'h2):(1'h1)]) ^~ (~^($unsigned(forvar916) ?
                      $unsigned(reg703) : reg892))) ?
                  (reg904[(3'h5):(2'h2)] >= (7'h47)) : (reg898[(4'h8):(1'h0)] & $unsigned($signed((reg765 < (8'hb0))))));
              reg924 <= reg686;
            end
        end
      reg925 = reg703[(3'h5):(1'h1)];
      if ({({reg741[(3'h4):(1'h1)]} ?
              $unsigned(((reg755 ?
                  reg715 : reg749) + (reg723 >> (8'hbc)))) : reg891[(4'ha):(1'h0)]),
          $unsigned(reg723[(3'h7):(3'h7)])})
        begin
          for (forvar926 = (1'h0); (forvar926 < (2'h2)); forvar926 = (forvar926 + (1'h1)))
            begin
              reg927 = reg771[(4'h8):(2'h3)];
              reg928 = $signed((reg739[(3'h5):(2'h2)] ?
                  (reg892[(3'h7):(3'h5)] != $unsigned(reg927)) : wire681));
            end
          if ((~|((reg928 ?
                  $unsigned((&reg696)) : $signed((reg898 && reg691))) ?
              reg697 : reg701[(3'h4):(3'h4)])))
            begin
              reg929 = $signed(reg920[(5'h13):(3'h6)]);
              reg930 <= $unsigned(((|($signed(reg922) != (~reg686))) < wire681));
              reg931 <= (($unsigned({{reg749}}) ?
                  {$unsigned($unsigned(reg899))} : {$signed((reg905 ?
                          reg924 : reg737)),
                      (8'hb8)}) != $signed((8'h9d)));
            end
          else
            begin
              reg930 <= $signed(reg708);
            end
          reg932 <= ($signed((~&$signed(((8'ha3) << (8'had))))) ?
              ($unsigned(reg739[(3'h4):(2'h3)]) & (~(~&$unsigned(reg888)))) : reg693[(3'h7):(2'h3)]);
          reg933 <= $unsigned(reg771[(1'h1):(1'h1)]);
        end
      else
        begin
          reg926 = reg880[(5'h11):(3'h7)];
          for (forvar927 = (1'h0); (forvar927 < (2'h3)); forvar927 = (forvar927 + (1'h1)))
            begin
              reg928 = reg737[(2'h3):(1'h1)];
              reg930 <= (reg920[(3'h7):(1'h0)] ?
                  $unsigned($signed(($signed(reg919) > wire872))) : (~&$signed((reg908 | reg743[(1'h1):(1'h0)]))));
              reg934 = wire680[(1'h1):(1'h0)];
              reg935 <= reg722[(4'ha):(2'h2)];
            end
          reg936 <= $unsigned(($unsigned($unsigned(reg919)) >= reg927[(1'h1):(1'h0)]));
        end
    end
  module937 #() modinst1139 (.wire939(reg702), .clk(clk), .y(wire1138), .wire940(reg707), .wire941(reg898), .wire938(reg722));
  always
    @(posedge clk) begin
      reg1140 <= reg936[(3'h6):(2'h3)];
      reg1141 <= ((^reg694[(4'h9):(3'h4)]) < (~(reg914[(4'hb):(3'h5)] ?
          reg904 : $unsigned($unsigned(reg737)))));
    end
  module1142 #() modinst1336 (.wire1145(reg691), .wire1146(reg703), .clk(clk), .y(wire1335), .wire1144(reg772), .wire1143(reg905), .wire1147(reg747));
  assign wire1337 = $unsigned(((~^($unsigned(reg697) ?
                        wire680[(1'h0):(1'h0)] : (reg707 ?
                            reg931 : reg932))) >>> (!reg931)));
  always
    @(posedge clk) begin
      reg1338 <= (reg746 >= (!((reg688[(2'h2):(1'h1)] ~^ {reg704}) >> {(+reg922)})));
      reg1339 = (~&reg924[(4'ha):(3'h4)]);
      for (forvar1340 = (1'h0); (forvar1340 < (1'h0)); forvar1340 = (forvar1340 + (1'h1)))
        begin
          for (forvar1341 = (1'h0); (forvar1341 < (2'h3)); forvar1341 = (forvar1341 + (1'h1)))
            begin
              reg1342 = $unsigned(((reg924[(2'h3):(1'h1)] + (&reg883)) ~^ (&((reg696 < reg749) != reg765))));
            end
        end
      reg1343 = reg755[(3'h7):(3'h5)];
      reg1344 = (~|reg740[(5'h12):(3'h5)]);
    end
  always
    @(posedge clk) begin
      reg1345 <= (reg920 ^~ ($signed($unsigned({(8'had), reg748})) ?
          (((wire1335 ? reg1140 : reg892) - $signed(reg907)) != (^(reg686 ?
              (8'ha4) : reg918))) : (($signed(reg712) ?
                  $unsigned(reg879) : (reg722 ? reg755 : reg722)) ?
              $unsigned({reg701, reg918}) : ($unsigned((8'hb7)) ?
                  reg734 : (8'h9f)))));
      reg1346 = (((reg694[(3'h4):(1'h0)] && {reg1338}) ^ reg743[(4'h9):(2'h3)]) ?
          wire1335 : (&reg935));
    end
  always
    @(posedge clk) begin
      reg1347 = $unsigned($unsigned(reg876[(1'h0):(1'h0)]));
      reg1348 = reg933;
      reg1349 <= {$unsigned($unsigned($signed((reg748 ? (8'hb9) : reg727)))),
          wire1335[(5'h10):(2'h2)]};
      reg1350 <= $unsigned(reg918[(1'h0):(1'h0)]);
      if ($signed($signed($unsigned((reg723 * $unsigned(reg697))))))
        begin
          reg1351 <= wire683[(5'h13):(4'hd)];
        end
      else
        begin
          reg1351 <= (^~(~$unsigned($signed($signed(wire680)))));
          for (forvar1352 = (1'h0); (forvar1352 < (1'h0)); forvar1352 = (forvar1352 + (1'h1)))
            begin
              reg1353 <= (wire684 ?
                  (~&(-(reg740[(1'h1):(1'h0)] >> (^~reg922)))) : ((reg702[(4'he):(2'h3)] == ({reg704,
                      reg922} >>> $signed(reg697))) >>> reg746));
              reg1354 = $signed($unsigned(reg1338));
              reg1355 <= (^((((~^reg922) << $unsigned(reg1350)) ?
                      ($unsigned(reg1345) ? {(8'hb2)} : (8'hb4)) : reg1350) ?
                  (reg891[(4'ha):(2'h3)] ?
                      ((reg902 >= wire683) < $unsigned(reg898)) : ((reg933 ?
                          reg718 : reg734) >> $unsigned((8'h9c)))) : (((|reg702) + (~|reg696)) ?
                      $signed({reg727}) : reg755[(3'h4):(2'h3)])));
              reg1356 = (~&{$unsigned((8'hb8))});
            end
          for (forvar1357 = (1'h0); (forvar1357 < (3'h4)); forvar1357 = (forvar1357 + (1'h1)))
            begin
              reg1358 <= $unsigned((reg718[(4'hb):(3'h5)] ?
                  {(8'hb5), reg704} : (~&$unsigned(reg708[(3'h7):(1'h1)]))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1359 = (1'h0); (forvar1359 < (1'h1)); forvar1359 = (forvar1359 + (1'h1)))
        begin
          for (forvar1360 = (1'h0); (forvar1360 < (2'h2)); forvar1360 = (forvar1360 + (1'h1)))
            begin
              reg1361 <= $unsigned($signed($signed(((reg712 ?
                  reg914 : wire1335) >>> reg1355))));
              reg1362 <= (&$unsigned((reg722 ?
                  {reg730, $unsigned(reg688)} : $signed($unsigned(wire682)))));
              reg1363 <= (((((8'hb0) ^ $unsigned(reg1350)) ?
                  {reg887} : reg876) || ($unsigned(reg686[(2'h3):(1'h0)]) ?
                  $signed(((7'h43) - reg740)) : {(reg924 ?
                          reg725 : reg712)})) > ((!reg887) ?
                  (-($unsigned(reg715) >>> reg712)) : reg932));
              reg1364 <= reg708[(3'h4):(1'h0)];
              reg1365 <= (^(reg1338[(1'h0):(1'h0)] > (((8'ha7) ^~ (^~reg755)) ?
                  reg1140 : reg1141)));
            end
          for (forvar1366 = (1'h0); (forvar1366 < (1'h1)); forvar1366 = (forvar1366 + (1'h1)))
            begin
              reg1367 = (~&$unsigned((!((forvar1360 ? (8'hbd) : reg876) ?
                  wire1138 : wire682))));
              reg1368 <= reg918[(3'h6):(3'h6)];
            end
          for (forvar1369 = (1'h0); (forvar1369 < (2'h2)); forvar1369 = (forvar1369 + (1'h1)))
            begin
              reg1370 <= (^~$signed($signed(((reg701 ~^ reg1361) <= $signed(reg688)))));
              reg1371 <= (~^$signed((reg898[(3'h4):(2'h2)] ~^ (reg923 ?
                  ((8'hb7) != reg1367) : (8'hbc)))));
            end
          for (forvar1372 = (1'h0); (forvar1372 < (1'h1)); forvar1372 = (forvar1372 + (1'h1)))
            begin
              reg1373 <= {reg734};
              reg1374 <= ($unsigned($signed((+((8'h9d) ? reg697 : reg887)))) ?
                  reg936[(4'hb):(4'h9)] : $signed(reg919));
              reg1375 = ({(~|reg703)} - reg930[(3'h7):(3'h4)]);
            end
          reg1376 <= ((^$unsigned(($signed(reg746) ?
                  $signed((8'ha7)) : (-reg1351)))) ?
              reg1358[(4'hd):(1'h0)] : (~&($unsigned($signed(reg730)) + reg1374)));
        end
      reg1377 = wire684[(4'hf):(2'h3)];
      reg1378 = (~^(+reg1355));
      for (forvar1379 = (1'h0); (forvar1379 < (3'h4)); forvar1379 = (forvar1379 + (1'h1)))
        begin
          reg1380 <= $unsigned({$unsigned($unsigned(wire683[(4'he):(4'h9)]))});
        end
    end
  always
    @(posedge clk) begin
      if ($signed(reg919[(3'h4):(3'h4)]))
        begin
          reg1381 <= $signed(($signed($signed({reg697})) ?
              (reg703[(4'hc):(4'hc)] ?
                  $signed($unsigned(wire872)) : (reg907[(3'h7):(3'h4)] + reg723[(4'h9):(4'h8)])) : reg924[(3'h4):(1'h0)]));
          for (forvar1382 = (1'h0); (forvar1382 < (1'h0)); forvar1382 = (forvar1382 + (1'h1)))
            begin
              reg1383 = reg1364;
              reg1384 = $signed(($unsigned(wire680[(4'hb):(4'h9)]) ?
                  $unsigned(reg887[(4'ha):(1'h0)]) : $signed(reg883[(2'h2):(1'h0)])));
            end
          for (forvar1385 = (1'h0); (forvar1385 < (1'h0)); forvar1385 = (forvar1385 + (1'h1)))
            begin
              reg1386 <= $signed(reg1384[(3'h7):(1'h1)]);
              reg1387 = ($signed((|reg1338[(1'h0):(1'h0)])) ?
                  (^~$signed(($unsigned(reg1351) ?
                      (^(8'hba)) : (reg686 << reg747)))) : reg1349);
            end
          if (reg1141[(3'h6):(3'h4)])
            begin
              reg1388 <= {$signed((reg708[(4'hc):(4'hc)] ?
                      $signed((~reg701)) : reg923[(3'h4):(2'h2)]))};
              reg1389 = reg722;
            end
          else
            begin
              reg1388 <= wire682;
              reg1390 <= ((((wire682[(3'h5):(3'h5)] - $unsigned((8'hac))) ^ (~(reg922 >= reg772))) | $unsigned(((reg1353 & reg688) << $unsigned(reg1383)))) ~^ ((-{(wire680 | wire1335),
                  ((8'hb0) ^~ reg1364)}) << $signed((reg771 & $unsigned(reg691)))));
            end
          for (forvar1391 = (1'h0); (forvar1391 < (1'h0)); forvar1391 = (forvar1391 + (1'h1)))
            begin
              reg1392 <= (~^$unsigned({($signed(reg1355) ?
                      $unsigned((7'h43)) : $signed(reg772))}));
              reg1393 <= reg737;
              reg1394 <= (reg1361[(1'h1):(1'h0)] | ((($signed(reg718) ?
                          (~&reg723) : reg883[(3'h4):(1'h1)]) ?
                      {reg883} : ((reg1390 ? (8'ha9) : reg1384) ?
                          (8'hb2) : (reg701 * reg734))) ?
                  (~^$unsigned({reg922})) : (~^$unsigned((reg898 ^ wire683)))));
            end
        end
      else
        begin
          reg1382 = reg1376;
        end
      if ((8'hb5))
        begin
          reg1395 = $unsigned({reg923[(2'h2):(1'h1)]});
          for (forvar1396 = (1'h0); (forvar1396 < (1'h0)); forvar1396 = (forvar1396 + (1'h1)))
            begin
              reg1397 <= (!(~|((-(reg772 ?
                  reg712 : reg725)) <<< $unsigned((wire684 ?
                  reg932 : reg694)))));
              reg1398 <= (&$signed((wire683[(3'h7):(3'h4)] != $unsigned((+reg1345)))));
              reg1399 = reg936[(2'h3):(1'h1)];
            end
          for (forvar1400 = (1'h0); (forvar1400 < (3'h4)); forvar1400 = (forvar1400 + (1'h1)))
            begin
              reg1401 <= ((reg1345 >= (reg1368 ?
                  $signed(((8'hb4) ?
                      (8'haa) : reg708)) : reg693[(2'h3):(1'h0)])) ^ (+{$unsigned(reg691)}));
            end
          if ($unsigned((+reg902[(4'h8):(1'h0)])))
            begin
              reg1402 <= $unsigned(((8'ha9) * (-$signed(reg908[(3'h4):(3'h4)]))));
              reg1403 = (|$unsigned(((~^$unsigned(reg1383)) != reg734)));
              reg1404 = (reg922 <<< (~^$signed((~&(wire683 - reg1345)))));
              reg1405 <= $unsigned(reg1404[(1'h1):(1'h0)]);
              reg1406 = {($unsigned($unsigned(wire1138[(4'hb):(3'h7)])) ?
                      ($signed((reg1374 ? reg691 : reg707)) ?
                          $signed($unsigned(reg935)) : $signed((reg899 < reg920))) : reg1349[(4'h8):(1'h0)]),
                  (reg898 + reg730)};
            end
          else
            begin
              reg1402 <= (~|$signed((+(|(~|(8'hb4))))));
              reg1405 <= reg747[(4'hd):(4'hc)];
              reg1407 <= $signed(reg701[(5'h14):(3'h4)]);
              reg1408 <= {$signed(({reg876} > (~(reg1381 < reg879))))};
            end
          for (forvar1409 = (1'h0); (forvar1409 < (1'h1)); forvar1409 = (forvar1409 + (1'h1)))
            begin
              reg1410 = (~&(^~($unsigned((reg1353 ? reg748 : (8'ha7))) ?
                  ((8'ha8) + reg702) : (reg765[(3'h5):(2'h2)] * (^~reg708)))));
              reg1411 = reg1383[(4'ha):(1'h0)];
              reg1412 <= ((~|($unsigned($unsigned((8'ha0))) >>> ($unsigned(reg931) >>> {reg746}))) ?
                  reg1395 : (((((8'hb3) ? reg776 : reg1368) >= (reg721 ?
                              reg1361 : reg748)) ?
                          $unsigned((^reg1358)) : reg931[(4'h9):(1'h0)]) ?
                      $unsigned(reg931) : (|forvar1396[(3'h4):(1'h0)])));
            end
        end
      else
        begin
          if ($signed({$signed((~|{wire1138})),
              ((|reg723[(4'he):(4'he)]) ?
                  (|$signed(reg1408)) : ((reg1368 ? reg904 : reg740) ?
                      (wire683 != reg739) : $signed(reg1398)))}))
            begin
              reg1396 <= {$signed(reg1412)};
              reg1399 = $signed(reg704[(4'hc):(3'h7)]);
              reg1400 <= ($unsigned({(7'h42), reg739[(3'h6):(1'h0)]}) ?
                  $signed($signed(({reg1351,
                      (8'ha7)} >> $signed(reg905)))) : (reg1387[(2'h3):(1'h1)] <<< {reg1373}));
              reg1403 = (reg708 ?
                  (reg1410 << reg707[(4'hd):(2'h2)]) : (~^$unsigned(((~^reg703) & $unsigned(reg739)))));
              reg1404 = reg737;
            end
          else
            begin
              reg1395 = $signed({(~&$unsigned($signed(reg712))),
                  $unsigned($unsigned($unsigned((8'haf))))});
              reg1396 <= (reg1392 ~^ (reg1392[(1'h0):(1'h0)] ?
                  reg1361 : reg935));
              reg1397 <= $unsigned((reg691[(4'hb):(1'h1)] ?
                  (8'ha2) : $signed($signed($unsigned(wire681)))));
            end
          reg1406 = {forvar1396, reg748};
        end
      reg1413 <= ((reg930 ?
          $signed($signed(reg902)) : $unsigned(($unsigned(reg1376) ?
              $unsigned(reg1393) : reg688[(4'h8):(3'h6)]))) + (~reg1358[(2'h3):(2'h3)]));
      if ($unsigned({($unsigned($unsigned((8'h9f))) > $signed((reg686 ?
              (8'hb5) : reg1397)))}))
        begin
          for (forvar1414 = (1'h0); (forvar1414 < (1'h1)); forvar1414 = (forvar1414 + (1'h1)))
            begin
              reg1415 <= {$unsigned($unsigned(((forvar1409 || reg1392) ?
                      reg704[(4'h9):(4'h9)] : (~^reg1395)))),
                  {$unsigned((8'ha8))}};
              reg1416 <= $signed(reg923[(2'h2):(1'h0)]);
            end
          reg1417 <= ((-$signed(($signed(reg905) ?
              $unsigned(reg1353) : (reg922 || reg1141)))) >> {reg919[(4'ha):(4'h9)]});
          reg1418 <= {($unsigned((reg904 > $unsigned(reg1338))) == ((~|(8'h9d)) || (~|{reg933,
                  reg935})))};
        end
      else
        begin
          if ((~^((reg1395 ?
                  (-reg1408[(1'h1):(1'h1)]) : ((reg1397 ? reg704 : reg1365) ?
                      reg1403 : (forvar1385 ? forvar1409 : reg721))) ?
              $unsigned(reg1353) : $signed(reg1401[(1'h0):(1'h0)]))))
            begin
              reg1414 <= reg704;
              reg1415 <= $signed($signed((((reg1370 ?
                      reg755 : reg1388) <= (reg892 >>> reg920)) ?
                  (-reg772[(4'h8):(2'h3)]) : reg1400[(1'h1):(1'h1)])));
            end
          else
            begin
              reg1414 <= ($signed((7'h43)) <= $signed(reg1371[(4'h9):(1'h1)]));
              reg1419 = ((!(reg914 ?
                      ((~^(8'hbc)) ?
                          $unsigned(reg718) : reg1380[(5'h11):(4'hf)]) : (-$signed(reg1355)))) ?
                  ((reg1406[(4'h8):(4'h8)] != reg739[(3'h4):(1'h0)]) >>> (~&$signed({reg688,
                      reg1370}))) : (~|(~&(|$signed(reg1351)))));
            end
        end
      for (forvar1420 = (1'h0); (forvar1420 < (3'h4)); forvar1420 = (forvar1420 + (1'h1)))
        begin
          if (reg936[(1'h0):(1'h0)])
            begin
              reg1421 <= (~&($signed(reg1363) ?
                  (~^($unsigned(reg688) ?
                      (!reg924) : reg1394[(1'h0):(1'h0)])) : ((-(reg730 ?
                          reg1364 : reg697)) ?
                      reg1392[(3'h7):(2'h2)] : (-$unsigned(reg1411)))));
            end
          else
            begin
              reg1421 <= $signed(reg1345[(2'h3):(2'h3)]);
            end
          if ((~^((+(-(reg739 ?
              reg1358 : (7'h44)))) * (((reg741 ~^ reg1390) < reg923[(1'h1):(1'h1)]) || $signed($unsigned(reg697))))))
            begin
              reg1422 <= reg1140;
            end
          else
            begin
              reg1423 = {(((&reg887[(4'ha):(3'h5)]) ?
                          $signed(reg771[(4'hb):(2'h2)]) : (reg1383 >> reg1363)) ?
                      {reg1140} : (forvar1420 ?
                          (!reg765[(2'h3):(2'h3)]) : reg931)),
                  reg1383[(1'h1):(1'h1)]};
              reg1424 <= ($signed(forvar1391) ?
                  reg734[(4'h8):(1'h0)] : (~|((reg1397 << $signed(forvar1382)) >> $unsigned(reg707))));
            end
          for (forvar1425 = (1'h0); (forvar1425 < (1'h0)); forvar1425 = (forvar1425 + (1'h1)))
            begin
              reg1426 <= $signed(((({forvar1391, reg1424} ?
                          (^reg1410) : (reg936 & reg1141)) ?
                      (!reg899) : $unsigned(reg765[(4'hd):(4'h8)])) ?
                  reg902[(3'h5):(3'h4)] : $unsigned($unsigned(reg1361[(2'h3):(2'h2)]))));
              reg1427 <= (reg1392 ?
                  $unsigned($unsigned(((8'hb5) ?
                      (reg1426 ?
                          forvar1385 : reg743) : (reg746 ~^ (8'hb3))))) : {$unsigned($signed((reg883 & forvar1409)))});
              reg1428 <= reg721;
              reg1429 <= (^$signed({forvar1414}));
            end
          reg1430 <= reg749[(3'h6):(2'h2)];
        end
    end
  assign wire1431 = $signed(reg694[(1'h0):(1'h0)]);
  module1432 #() modinst1594 (wire1593, clk, reg902, reg718, reg1351, reg725);
  assign wire1595 = ($signed((&(((8'h9d) > reg725) ?
                            $signed(reg936) : (reg1376 ? reg1414 : reg694)))) ?
                        (!$unsigned(((~reg1368) & {reg1415}))) : $signed(reg1418[(1'h1):(1'h1)]));
  always
    @(posedge clk) begin
      reg1596 <= (reg1365 | reg1417[(3'h4):(2'h3)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module71  (y, clk, wire72, wire73, wire74, wire75);
  output wire [(32'h725):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire72;
  input wire signed [(4'hb):(1'h0)] wire73;
  input wire signed [(3'h6):(1'h0)] wire74;
  input wire signed [(5'h15):(1'h0)] wire75;
  wire [(3'h6):(1'h0)] wire658;
  wire [(3'h6):(1'h0)] wire657;
  wire [(4'hd):(1'h0)] wire656;
  wire signed [(5'h16):(1'h0)] wire654;
  wire [(5'h16):(1'h0)] wire521;
  wire [(3'h6):(1'h0)] wire76;
  wire signed [(5'h14):(1'h0)] wire77;
  wire [(4'hd):(1'h0)] wire78;
  wire signed [(2'h2):(1'h0)] wire94;
  wire [(5'h14):(1'h0)] wire140;
  wire signed [(3'h6):(1'h0)] wire508;
  reg signed [(5'h12):(1'h0)] reg187 = (1'h0);
  reg [(5'h13):(1'h0)] reg192 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg189 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg188 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg186 = (1'h0);
  reg [(4'hc):(1'h0)] reg183 = (1'h0);
  reg [(4'h9):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg180 = (1'h0);
  reg [(4'hd):(1'h0)] reg179 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg178 = (1'h0);
  reg [(3'h4):(1'h0)] reg177 = (1'h0);
  reg [(5'h14):(1'h0)] reg176 = (1'h0);
  reg [(5'h10):(1'h0)] reg175 = (1'h0);
  reg [(5'h17):(1'h0)] reg172 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg170 = (1'h0);
  reg [(5'h16):(1'h0)] reg169 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg156 = (1'h0);
  reg [(3'h5):(1'h0)] reg155 = (1'h0);
  reg [(5'h13):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg148 = (1'h0);
  reg [(5'h16):(1'h0)] reg147 = (1'h0);
  reg [(4'h9):(1'h0)] reg146 = (1'h0);
  reg [(4'he):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg144 = (1'h0);
  reg [(3'h7):(1'h0)] reg142 = (1'h0);
  reg [(3'h4):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg138 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg137 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg136 = (1'h0);
  reg [(5'h10):(1'h0)] reg134 = (1'h0);
  reg [(4'h8):(1'h0)] reg130 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg128 = (1'h0);
  reg [(4'hf):(1'h0)] reg125 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg124 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg122 = (1'h0);
  reg [(5'h15):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg119 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg116 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg109 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg108 = (1'h0);
  reg [(5'h10):(1'h0)] reg103 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg101 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg99 = (1'h0);
  reg [(5'h17):(1'h0)] reg98 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg97 = (1'h0);
  reg [(4'hd):(1'h0)] reg95 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg93 = (1'h0);
  reg [(2'h3):(1'h0)] reg92 = (1'h0);
  reg [(3'h4):(1'h0)] reg90 = (1'h0);
  reg [(5'h15):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg84 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg81 = (1'h0);
  reg [(2'h3):(1'h0)] reg79 = (1'h0);
  reg [(4'h8):(1'h0)] reg510 = (1'h0);
  reg [(4'hd):(1'h0)] reg511 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg512 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg514 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg515 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg517 = (1'h0);
  reg [(3'h4):(1'h0)] reg519 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg520 = (1'h0);
  reg [(5'h10):(1'h0)] forvar512 = (1'h0);
  reg [(5'h15):(1'h0)] reg518 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg516 = (1'h0);
  reg [(4'hf):(1'h0)] reg513 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg194 = (1'h0);
  reg [(4'hf):(1'h0)] forvar193 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg191 = (1'h0);
  reg [(5'h15):(1'h0)] reg190 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar187 = (1'h0);
  reg [(4'hc):(1'h0)] reg185 = (1'h0);
  reg [(3'h4):(1'h0)] reg184 = (1'h0);
  reg [(5'h13):(1'h0)] reg181 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg174 = (1'h0);
  reg signed [(4'he):(1'h0)] reg173 = (1'h0);
  reg [(5'h14):(1'h0)] forvar171 = (1'h0);
  reg [(5'h10):(1'h0)] reg168 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg167 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg166 = (1'h0);
  reg [(5'h14):(1'h0)] reg165 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar164 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar163 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg162 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar161 = (1'h0);
  reg [(2'h3):(1'h0)] reg160 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar159 = (1'h0);
  reg [(4'h9):(1'h0)] reg158 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar157 = (1'h0);
  reg signed [(4'he):(1'h0)] reg154 = (1'h0);
  reg [(3'h4):(1'h0)] reg152 = (1'h0);
  reg signed [(4'he):(1'h0)] reg151 = (1'h0);
  reg [(3'h4):(1'h0)] forvar150 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg149 = (1'h0);
  reg [(4'he):(1'h0)] reg143 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar141 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar135 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar133 = (1'h0);
  reg [(4'hf):(1'h0)] reg132 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg131 = (1'h0);
  reg [(5'h12):(1'h0)] reg129 = (1'h0);
  reg [(4'he):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg126 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar121 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar118 = (1'h0);
  reg [(4'hd):(1'h0)] reg117 = (1'h0);
  reg [(2'h2):(1'h0)] forvar115 = (1'h0);
  reg [(3'h4):(1'h0)] reg114 = (1'h0);
  reg [(5'h13):(1'h0)] reg113 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg112 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg111 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg107 = (1'h0);
  reg [(5'h13):(1'h0)] reg106 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg105 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg104 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg102 = (1'h0);
  reg [(4'he):(1'h0)] reg100 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar96 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg91 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg89 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg88 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg87 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg85 = (1'h0);
  reg [(5'h14):(1'h0)] forvar83 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg82 = (1'h0);
  reg [(5'h10):(1'h0)] forvar80 = (1'h0);
  assign y = {wire658,
                 wire657,
                 wire656,
                 wire654,
                 wire521,
                 wire76,
                 wire77,
                 wire78,
                 wire94,
                 wire140,
                 wire508,
                 reg187,
                 reg192,
                 reg189,
                 reg188,
                 reg186,
                 reg183,
                 reg182,
                 reg180,
                 reg179,
                 reg178,
                 reg177,
                 reg176,
                 reg175,
                 reg172,
                 reg170,
                 reg169,
                 reg156,
                 reg155,
                 reg153,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg142,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg134,
                 reg130,
                 reg128,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg120,
                 reg119,
                 reg116,
                 reg109,
                 reg108,
                 reg103,
                 reg101,
                 reg99,
                 reg98,
                 reg97,
                 reg95,
                 reg93,
                 reg92,
                 reg90,
                 reg86,
                 reg84,
                 reg81,
                 reg79,
                 reg510,
                 reg511,
                 reg512,
                 reg514,
                 reg515,
                 reg517,
                 reg519,
                 reg520,
                 forvar512,
                 reg518,
                 reg516,
                 reg513,
                 reg193,
                 reg194,
                 forvar193,
                 reg191,
                 reg190,
                 forvar187,
                 reg185,
                 reg184,
                 reg181,
                 reg174,
                 reg173,
                 forvar171,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 forvar164,
                 forvar163,
                 reg162,
                 forvar161,
                 reg160,
                 forvar159,
                 reg158,
                 forvar157,
                 reg154,
                 reg152,
                 reg151,
                 forvar150,
                 reg149,
                 reg143,
                 forvar141,
                 forvar135,
                 forvar133,
                 reg132,
                 reg131,
                 reg129,
                 reg127,
                 reg126,
                 forvar121,
                 forvar118,
                 reg117,
                 forvar115,
                 reg114,
                 reg113,
                 reg112,
                 reg111,
                 reg110,
                 reg107,
                 reg106,
                 reg105,
                 reg104,
                 reg102,
                 reg100,
                 forvar96,
                 reg91,
                 reg89,
                 reg88,
                 reg87,
                 reg85,
                 forvar83,
                 reg82,
                 forvar80,
                 (1'h0)};
  assign wire76 = (wire75 ?
                      (wire75 >>> ($signed($signed(wire72)) ?
                          (-(7'h47)) : $unsigned(((8'haf) ?
                              (8'hae) : wire73)))) : (wire74 ?
                          $signed((((8'h9f) ~^ (8'hbe)) + wire72)) : (8'h9e)));
  assign wire77 = (($unsigned($unsigned(wire73[(2'h2):(1'h1)])) > $signed(((wire74 == wire73) ?
                      $unsigned(wire76) : $unsigned(wire73)))) << wire76);
  assign wire78 = (8'hb4);
  always
    @(posedge clk) begin
      reg79 <= (~&($signed(wire75) ?
          (~(^(wire75 ? (8'hb8) : wire73))) : (~|wire77)));
      for (forvar80 = (1'h0); (forvar80 < (2'h3)); forvar80 = (forvar80 + (1'h1)))
        begin
          reg81 <= (~^((wire73 & ($signed(wire75) ?
              {(8'ha7)} : (wire72 ?
                  wire75 : (7'h48)))) + $unsigned((+wire78[(1'h0):(1'h0)]))));
          reg82 = $signed($signed(wire74[(2'h2):(1'h0)]));
          for (forvar83 = (1'h0); (forvar83 < (2'h3)); forvar83 = (forvar83 + (1'h1)))
            begin
              reg84 <= (&$signed({wire75[(3'h5):(2'h2)]}));
            end
          if ((~(reg82 ?
              {$signed($unsigned(reg82))} : (+$signed(((8'hb7) >> (7'h45)))))))
            begin
              reg85 = $signed({{{{reg82, reg84}},
                      ({forvar83, wire78} ?
                          wire74[(1'h0):(1'h0)] : (~(7'h4a)))}});
            end
          else
            begin
              reg85 = $unsigned(wire74);
              reg86 <= $signed(((~($unsigned(wire78) ?
                  reg79 : $signed(wire74))) ^ {$unsigned((~^wire72))}));
              reg87 = ((wire75 ?
                  $unsigned(reg81) : $unsigned($signed(reg81[(5'h16):(5'h13)]))) < wire74[(2'h3):(2'h3)]);
              reg88 = ({$signed({(~reg85), {(8'ha3), reg86}}),
                  (forvar80 ?
                      $signed($signed(wire73)) : $signed($unsigned(reg82)))} - wire77);
              reg89 = {(&(~^reg84)), reg86[(5'h13):(3'h5)]};
            end
          if ((forvar80[(4'he):(2'h3)] < $unsigned(wire75)))
            begin
              reg90 <= $signed((^($signed((~wire75)) ?
                  ($unsigned(reg86) ? (reg82 << wire75) : forvar83) : ({wire72,
                      wire78} != (~reg87)))));
            end
          else
            begin
              reg90 <= $unsigned({{reg79, forvar83}});
              reg91 = ((8'ha0) & (~&reg87));
              reg92 <= $unsigned(reg89);
              reg93 <= (((^~$unsigned($unsigned(wire76))) || wire72[(4'he):(1'h1)]) | (((wire78[(3'h5):(1'h1)] & wire75[(4'ha):(1'h0)]) <= ($signed(reg86) ?
                  wire78 : reg86)) ^ {(wire72 ?
                      (wire76 ^ reg81) : $unsigned(forvar83))}));
            end
        end
    end
  assign wire94 = (reg84[(4'h9):(3'h7)] & $signed($unsigned(reg81[(2'h2):(2'h2)])));
  always
    @(posedge clk) begin
      reg95 <= (~$unsigned(reg90));
      for (forvar96 = (1'h0); (forvar96 < (1'h0)); forvar96 = (forvar96 + (1'h1)))
        begin
          reg97 <= $unsigned($unsigned($unsigned($unsigned(wire94))));
          if ((^~$unsigned(({{wire94}} < $signed((reg79 ? wire94 : wire77))))))
            begin
              reg98 <= $unsigned(($signed((8'hb9)) ?
                  $signed($unsigned((wire77 | (8'hbf)))) : ((reg84[(2'h3):(1'h0)] ?
                          (^~wire94) : $signed(wire74)) ?
                      (~(^~wire72)) : {(8'hbd), $unsigned((8'ha0))})));
              reg99 <= (($signed({reg93[(5'h14):(4'hd)], {wire74, reg81}}) ?
                  $signed((~^$unsigned(wire73))) : (((wire73 ?
                          wire72 : reg84) || reg95[(3'h6):(3'h4)]) ?
                      (+reg86) : (8'hbe))) + ($unsigned(forvar96) ?
                  $signed(reg92[(1'h0):(1'h0)]) : ({(reg92 <<< wire74),
                          $unsigned(reg95)} ?
                      {wire76,
                          (wire77 ? reg98 : reg93)} : (+$unsigned(reg81)))));
              reg100 = $signed({reg97[(3'h6):(3'h6)], wire94});
              reg101 <= (reg86 ?
                  reg81[(4'h9):(1'h1)] : ($signed((reg100 <<< wire77)) ?
                      ((wire72 ?
                          $unsigned(reg92) : $signed(reg79)) << forvar96[(4'h9):(1'h1)]) : (|reg81)));
            end
          else
            begin
              reg98 <= wire74;
              reg100 = wire77[(4'hc):(4'hb)];
              reg102 = (($signed($unsigned(reg84)) * ((^(reg95 ^~ wire94)) < reg84)) == ($signed($unsigned((reg99 ~^ reg93))) + $unsigned({$unsigned(wire94),
                  {reg95, wire94}})));
            end
          reg103 <= $signed((reg97[(2'h2):(1'h1)] || {$unsigned(reg93),
              $signed($unsigned(reg101))}));
        end
      reg104 = wire76;
      if ((-reg100))
        begin
          if (reg93[(4'hd):(4'hd)])
            begin
              reg105 = $signed((reg86[(3'h4):(2'h3)] || (|((wire94 ?
                  wire94 : wire72) != reg79))));
              reg106 = $signed(reg93[(5'h12):(5'h12)]);
              reg107 = $unsigned($unsigned(reg101[(3'h5):(2'h3)]));
            end
          else
            begin
              reg105 = ((+reg103[(4'hf):(3'h7)]) ?
                  reg90[(1'h0):(1'h0)] : $signed($signed(($signed(reg97) ?
                      (&reg104) : (-reg103)))));
              reg106 = {(^wire78[(4'hb):(3'h6)]), (~^reg93[(4'ha):(4'ha)])};
              reg108 <= $unsigned($signed((reg93[(5'h16):(4'hb)] ?
                  (((8'ha6) ? reg81 : reg103) || {reg107}) : (+(reg90 ?
                      (8'ha0) : reg92)))));
              reg109 <= $signed((reg106 ?
                  (((!reg105) ? $signed(reg79) : (~|forvar96)) ?
                      ($unsigned((7'h45)) < wire72[(3'h4):(1'h1)]) : wire94[(2'h2):(2'h2)]) : $signed($signed(reg107))));
            end
          reg110 = wire72;
          if ((((8'ha9) ?
                  $signed({(7'h43)}) : {(forvar96 + (&(7'h49))),
                      ($signed(wire72) ? {reg95} : (wire73 ? reg92 : reg98))}) ?
              reg99 : $unsigned($unsigned({(reg86 ~^ wire74), reg103}))))
            begin
              reg111 = (reg105 >> $unsigned($unsigned(((8'ha8) + (+reg107)))));
              reg112 = $unsigned($signed((~$signed((8'ha4)))));
              reg113 = (reg111[(2'h3):(2'h3)] ?
                  reg112 : ($unsigned((~|(forvar96 ?
                      (8'hab) : reg101))) ^~ ({(~&reg107),
                          wire78[(4'ha):(3'h7)]} ?
                      $unsigned((reg99 ?
                          wire94 : reg100)) : $unsigned(reg86))));
              reg114 = {((($signed(reg113) ? $unsigned(wire72) : (7'h49)) ?
                      $signed((~^wire73)) : ($unsigned(wire76) != (reg106 >> reg79))) != (|reg112)),
                  $unsigned((&((~|wire94) ?
                      $unsigned((8'ha8)) : reg81[(4'hf):(4'he)])))};
            end
          else
            begin
              reg111 = (+reg104[(1'h1):(1'h0)]);
              reg112 = reg109[(5'h10):(4'he)];
              reg113 = (($unsigned((reg114[(2'h2):(1'h0)] ~^ reg107)) ?
                      $signed($unsigned((-reg107))) : $signed(((^reg112) <<< (reg79 ?
                          wire77 : reg98)))) ?
                  {{(&wire94)}, (&reg114)} : wire78);
            end
        end
      else
        begin
          reg105 = reg84;
          reg108 <= reg93[(4'hc):(4'hc)];
          reg109 <= (reg109 ?
              (reg95[(3'h4):(3'h4)] && $signed($unsigned(wire77))) : reg98[(5'h10):(3'h4)]);
        end
      for (forvar115 = (1'h0); (forvar115 < (2'h2)); forvar115 = (forvar115 + (1'h1)))
        begin
          reg116 <= $signed($signed((~^$signed((+reg103)))));
        end
    end
  always
    @(posedge clk) begin
      reg117 = (+((~^$signed((reg103 ? reg109 : reg86))) ?
          $unsigned($signed(reg108[(1'h0):(1'h0)])) : reg93[(4'hd):(1'h0)]));
    end
  always
    @(posedge clk) begin
      for (forvar118 = (1'h0); (forvar118 < (2'h3)); forvar118 = (forvar118 + (1'h1)))
        begin
          reg119 <= $signed($signed($unsigned((-(&(8'hac))))));
          reg120 <= ((reg97 ?
              ({$unsigned((7'h4a)),
                  (~^reg79)} > $signed($unsigned((8'hb4)))) : ((^((8'hb6) ?
                  reg116 : reg81)) ~^ ((^wire75) ?
                  $signed(reg99) : $unsigned(wire73)))) != wire72[(5'h14):(4'he)]);
          for (forvar121 = (1'h0); (forvar121 < (2'h2)); forvar121 = (forvar121 + (1'h1)))
            begin
              reg122 <= (!$signed($unsigned(((reg79 ?
                  reg86 : reg92) ~^ $signed(wire78)))));
            end
          if ((^~(~(~{wire94}))))
            begin
              reg123 <= {forvar121, reg95};
              reg124 <= reg120;
              reg125 <= ((~|reg101) <<< ((8'h9f) <= $signed(wire76)));
            end
          else
            begin
              reg126 = wire73[(1'h1):(1'h1)];
            end
          if ($unsigned(reg103[(4'hd):(4'hc)]))
            begin
              reg127 = reg109[(1'h1):(1'h1)];
              reg128 <= $signed(wire77[(4'hf):(3'h5)]);
              reg129 = $signed(($signed($unsigned((reg99 ~^ reg125))) ~^ (~$unsigned((wire76 != reg86)))));
              reg130 <= $signed((8'ha9));
            end
          else
            begin
              reg127 = ((((-forvar121[(2'h3):(1'h0)]) != (8'ha1)) ?
                      reg92[(2'h2):(1'h0)] : (8'h9d)) ?
                  (^~reg119) : $unsigned((reg95[(3'h5):(1'h0)] - wire75)));
              reg129 = forvar121;
              reg131 = {(&wire74)};
              reg132 = reg93;
            end
        end
      for (forvar133 = (1'h0); (forvar133 < (1'h0)); forvar133 = (forvar133 + (1'h1)))
        begin
          reg134 <= ($signed($unsigned(reg98)) ?
              (reg129[(2'h2):(2'h2)] || ($signed((wire94 ? reg97 : reg86)) ?
                  $signed(forvar133) : (((8'hae) ?
                      reg84 : reg97) ~^ ((8'haa) & forvar121)))) : ($unsigned($unsigned(reg90[(1'h0):(1'h0)])) ?
                  (reg125[(3'h7):(2'h2)] ?
                      (^~(8'ha6)) : $unsigned((reg125 ?
                          reg122 : reg132))) : (((+reg97) | (^(8'ha0))) ?
                      ((&reg109) ?
                          reg116[(4'hb):(3'h6)] : (~|reg95)) : ($signed(wire94) ?
                          $unsigned(reg122) : (~(8'had))))));
          for (forvar135 = (1'h0); (forvar135 < (3'h4)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 <= $signed(((wire77[(5'h12):(4'hb)] ?
                      $unsigned($signed(wire77)) : reg127[(2'h2):(1'h0)]) ?
                  {$unsigned(reg125[(3'h6):(1'h0)]),
                      $signed((8'hb0))} : reg103[(5'h10):(3'h6)]));
              reg137 <= (($signed(wire78) ? $unsigned(reg98) : reg124) ?
                  (({reg95, (^forvar135)} >> $unsigned($signed(reg127))) ?
                      reg108 : reg136[(4'h9):(2'h2)]) : $unsigned(reg90));
              reg138 <= ($unsigned({$signed(wire77), {$signed(reg99)}}) ?
                  ($unsigned((~|(wire75 >>> reg130))) & (^~reg92)) : (reg122 - (({reg101} ?
                      (wire75 ?
                          forvar121 : reg109) : reg99) && reg92[(1'h1):(1'h0)])));
            end
          reg139 <= $unsigned($unsigned($unsigned($unsigned((~(8'ha2))))));
        end
    end
  assign wire140 = reg79;
  always
    @(posedge clk) begin
      for (forvar141 = (1'h0); (forvar141 < (3'h4)); forvar141 = (forvar141 + (1'h1)))
        begin
          if (reg108[(3'h5):(3'h4)])
            begin
              reg142 <= {({$signed(wire74),
                          (wire73 ?
                              (reg90 ? reg130 : wire74) : (reg139 ?
                                  reg130 : reg93))} ?
                      reg139 : $signed(wire77)),
                  (((8'ha4) ?
                          ($signed(reg95) ?
                              ((8'hbd) ? reg109 : reg137) : (reg109 ?
                                  reg90 : wire78)) : ((reg99 ? wire76 : reg95) ?
                              (^~wire94) : reg103[(1'h0):(1'h0)])) ?
                      $signed(({reg122,
                          (8'had)} == {(8'had)})) : {{(forvar141 - (7'h47))},
                          reg101[(4'ha):(3'h7)]})};
              reg143 = (~&wire76[(3'h5):(2'h3)]);
              reg144 <= reg137[(3'h4):(1'h1)];
              reg145 <= wire75[(4'h8):(2'h3)];
            end
          else
            begin
              reg143 = $unsigned($signed($unsigned(reg144[(4'h8):(2'h2)])));
              reg144 <= reg144;
              reg145 <= {(8'ha2)};
            end
          if (((-reg125[(4'h9):(3'h7)]) ? $signed(reg101) : wire140))
            begin
              reg146 <= $signed($unsigned(((+$unsigned(reg143)) ?
                  reg139 : $signed($unsigned(reg136)))));
            end
          else
            begin
              reg146 <= {($signed($unsigned($unsigned(reg137))) && reg79),
                  reg145};
              reg147 <= (reg84[(3'h4):(3'h4)] ? reg97 : reg79[(2'h2):(1'h1)]);
            end
          reg148 <= $signed((8'haf));
          reg149 = (^~$unsigned($signed((+$signed((8'hb1))))));
          for (forvar150 = (1'h0); (forvar150 < (3'h4)); forvar150 = (forvar150 + (1'h1)))
            begin
              reg151 = (^{reg81[(4'he):(4'ha)],
                  (+{((7'h45) < reg137), $signed((8'hbd))})});
              reg152 = (~$signed((|{(reg116 > (7'h42))})));
              reg153 <= (^~reg134[(3'h6):(1'h0)]);
              reg154 = (^$signed(($unsigned($unsigned(reg137)) ?
                  $unsigned((reg92 <= reg120)) : $signed(reg134[(4'ha):(3'h4)]))));
              reg155 <= {$signed($unsigned($unsigned((&reg138))))};
            end
        end
      reg156 <= reg108;
      for (forvar157 = (1'h0); (forvar157 < (1'h1)); forvar157 = (forvar157 + (1'h1)))
        begin
          reg158 = reg149[(1'h1):(1'h0)];
          for (forvar159 = (1'h0); (forvar159 < (1'h0)); forvar159 = (forvar159 + (1'h1)))
            begin
              reg160 = $unsigned($signed((^~((wire72 ? reg120 : reg158) ?
                  (-reg142) : (&reg116)))));
            end
        end
      for (forvar161 = (1'h0); (forvar161 < (1'h0)); forvar161 = (forvar161 + (1'h1)))
        begin
          reg162 = (((8'ha7) ?
                  (~|$unsigned(reg145)) : (+((reg128 ? reg92 : reg92) ?
                      (~&reg158) : (wire74 ? (7'h4a) : reg119)))) ?
              (($signed((reg95 ? reg151 : reg122)) ?
                      (8'hb9) : {reg86, reg142[(3'h6):(1'h1)]}) ?
                  $unsigned((7'h48)) : (&reg143[(3'h6):(3'h6)])) : {$unsigned($unsigned((~^reg84))),
                  (~&$signed(reg137))});
        end
      for (forvar163 = (1'h0); (forvar163 < (3'h4)); forvar163 = (forvar163 + (1'h1)))
        begin
          for (forvar164 = (1'h0); (forvar164 < (3'h4)); forvar164 = (forvar164 + (1'h1)))
            begin
              reg165 = {$signed({((reg98 ? wire78 : wire76) ?
                          wire94 : (reg119 || forvar141))})};
              reg166 = {((+$unsigned((reg122 - (7'h42)))) ?
                      reg98[(5'h14):(3'h7)] : (($unsigned(wire74) ?
                              (reg155 * reg103) : $unsigned(reg98)) ?
                          reg84[(4'h8):(2'h3)] : ({reg139, reg95} ?
                              $unsigned(reg109) : forvar163))),
                  $signed(((^reg148) >>> ((-wire78) ?
                      $unsigned((8'hac)) : reg144[(4'h9):(3'h7)])))};
              reg167 = forvar157;
              reg168 = reg145[(4'h9):(3'h5)];
              reg169 <= (-(reg165[(5'h12):(2'h3)] ?
                  $signed(((~|forvar157) <<< reg166)) : reg149[(2'h3):(2'h3)]));
            end
          reg170 <= (reg120 | ((!wire77[(3'h5):(2'h3)]) ?
              $signed((~^reg103)) : $signed(((reg97 + reg146) >= (reg149 <= wire77)))));
          for (forvar171 = (1'h0); (forvar171 < (2'h3)); forvar171 = (forvar171 + (1'h1)))
            begin
              reg172 <= (forvar159 * reg167[(3'h5):(1'h0)]);
              reg173 = (($signed(((reg169 ? (8'ha4) : (7'h47)) - (wire94 ?
                      reg101 : reg138))) ?
                  $unsigned(($unsigned(reg116) || {reg146})) : reg123) != ({($signed(reg154) < $unsigned((8'h9e))),
                      reg153} ?
                  reg158[(4'h8):(3'h5)] : reg142));
            end
          reg174 = (({{(~|reg172), reg84[(3'h4):(2'h3)]},
              ({reg142, reg98} ?
                  {reg169,
                      forvar141} : (8'hb9))} == $unsigned($signed($signed(reg149)))) < reg160);
        end
    end
  always
    @(posedge clk) begin
      reg175 <= (((((reg95 + (8'hb9)) ? (reg116 < reg103) : wire78) ?
              $signed((reg81 >>> (8'ha5))) : (~|$unsigned(reg120))) & ((~|{reg123,
                  (7'h49)}) ?
              (((8'hba) ?
                  reg136 : reg125) >= $unsigned(reg101)) : $signed($unsigned(wire77)))) ?
          {$signed($unsigned((wire94 + reg84))),
              $signed(reg123[(2'h2):(2'h2)])} : ((|(|reg145)) ?
              ($unsigned((reg95 ?
                  reg156 : reg134)) | $signed(wire94)) : reg142[(3'h4):(2'h3)]));
      if ((|$unsigned((^$unsigned((reg97 ? reg99 : (8'ha4)))))))
        begin
          reg176 <= {(reg156[(3'h7):(2'h2)] > ((reg84 ?
                  (reg86 < reg146) : (|reg138)) >>> wire73))};
        end
      else
        begin
          reg176 <= (8'h9c);
          reg177 <= wire72[(4'he):(2'h2)];
          if ((((wire75 ^~ $unsigned((reg124 ? reg116 : reg93))) ?
              reg108[(3'h6):(1'h0)] : (reg120[(3'h7):(3'h6)] ?
                  {reg128[(1'h0):(1'h0)],
                      (+reg169)} : $signed($signed(reg101)))) || ($signed(($signed(wire78) ?
              (^~reg175) : reg130[(2'h3):(1'h0)])) < $unsigned((reg81 & (wire77 - wire94))))))
            begin
              reg178 <= $unsigned($signed((($signed(reg177) == reg176) ?
                  (|$signed(wire78)) : wire73[(3'h4):(1'h0)])));
            end
          else
            begin
              reg178 <= reg136;
              reg179 <= reg139[(2'h3):(1'h1)];
              reg180 <= (reg177[(2'h2):(1'h0)] - reg178[(3'h5):(2'h3)]);
              reg181 = (^~(reg138 == $unsigned(reg178[(2'h2):(1'h0)])));
            end
        end
      if ($unsigned(reg170))
        begin
          if (reg81[(5'h15):(1'h1)])
            begin
              reg182 <= reg177[(3'h4):(2'h2)];
              reg183 <= reg179;
              reg184 = $signed(($unsigned($signed(reg108[(4'h9):(3'h7)])) ?
                  $unsigned(($signed(reg181) ?
                      $signed(reg81) : wire74)) : $signed({$unsigned(reg170),
                      (|(8'ha8))})));
              reg185 = $unsigned($signed(reg128));
            end
          else
            begin
              reg184 = $signed(wire75);
              reg185 = $signed($signed($unsigned($unsigned($unsigned(reg153)))));
              reg186 <= $signed($unsigned($unsigned(((8'hb2) & $signed(reg84)))));
            end
          for (forvar187 = (1'h0); (forvar187 < (1'h0)); forvar187 = (forvar187 + (1'h1)))
            begin
              reg188 <= (^wire72[(5'h13):(5'h12)]);
              reg189 <= (~|(~&($unsigned($signed(reg179)) >>> wire73[(4'h8):(3'h5)])));
              reg190 = wire76[(2'h3):(2'h3)];
            end
          reg191 = ({{(&{reg103, reg109})}} || reg144[(2'h2):(1'h0)]);
          reg192 <= (|($unsigned(reg184[(1'h0):(1'h0)]) >>> wire74[(2'h2):(1'h0)]));
          for (forvar193 = (1'h0); (forvar193 < (3'h4)); forvar193 = (forvar193 + (1'h1)))
            begin
              reg194 = (&$unsigned($unsigned($signed($unsigned(wire74)))));
            end
        end
      else
        begin
          if (reg189[(2'h2):(1'h0)])
            begin
              reg182 <= (reg120[(3'h5):(1'h1)] >> (((((8'haf) ?
                          wire74 : reg139) ?
                      (reg136 >> wire72) : (reg179 <<< reg194)) ?
                  reg124 : (-{reg124})) >= wire77[(3'h4):(2'h3)]));
              reg184 = {$unsigned((+(((8'hb7) ?
                      wire76 : reg130) << {reg175})))};
              reg185 = ((~^((reg103[(2'h3):(1'h1)] ~^ reg98) ?
                  (~^$unsigned((8'hae))) : (8'hb1))) + (+$unsigned((~|reg139))));
            end
          else
            begin
              reg182 <= $signed({wire140[(3'h4):(1'h1)], reg124});
              reg183 <= $unsigned(reg130);
              reg184 = reg179[(1'h1):(1'h1)];
              reg186 <= (reg124[(2'h3):(1'h1)] - ({(reg90 ?
                      reg181[(5'h10):(4'ha)] : (reg190 - reg124)),
                  $signed((reg84 ^~ reg156))} ^~ {reg175}));
            end
          if (reg146)
            begin
              reg187 <= {reg109,
                  (|$signed(($signed(reg148) ? {wire140} : $signed(reg177))))};
            end
          else
            begin
              reg190 = ($unsigned(($signed((~|(8'h9d))) >> $unsigned((reg146 <= reg130)))) ?
                  (reg90 ^~ {((!reg189) ^ reg169[(4'ha):(1'h1)]),
                      reg136}) : $signed(reg175));
              reg192 <= reg186;
              reg193 = $unsigned(reg178[(1'h0):(1'h0)]);
            end
        end
    end
  module195 #() modinst509 (wire508, clk, reg109, reg86, wire75, reg153);
  always
    @(posedge clk) begin
      reg510 <= $unsigned($unsigned(reg108));
    end
  always
    @(posedge clk) begin
      reg511 <= ((!(~^wire94[(2'h2):(1'h0)])) ^~ $signed($unsigned(((!reg183) ^ reg81[(3'h7):(3'h5)]))));
      if ({{$unsigned($signed(reg187)), (8'haa)}})
        begin
          reg512 <= reg189;
          if (reg142[(3'h7):(1'h0)])
            begin
              reg513 = ($signed($unsigned((!(8'h9d)))) ?
                  $unsigned($unsigned((^reg179))) : ((|(^reg182)) || (((reg122 ?
                          reg144 : reg511) ?
                      (7'h4a) : $unsigned(wire140)) <= reg119[(1'h1):(1'h0)])));
              reg514 <= $signed((~|($unsigned((!reg172)) >= ($signed(reg95) + wire94))));
              reg515 <= reg155;
            end
          else
            begin
              reg513 = (-$signed($signed(((reg130 & (7'h48)) >= $unsigned(reg146)))));
              reg514 <= reg97[(4'h8):(3'h6)];
              reg515 <= ($unsigned((((reg188 ? (8'hbb) : reg514) < {reg182}) ?
                      $signed((reg124 ?
                          reg120 : wire78)) : reg148[(4'hd):(4'hb)])) ?
                  $unsigned((8'hb5)) : (reg179 ?
                      (+$unsigned((reg169 || reg180))) : reg95));
              reg516 = $unsigned(reg119[(4'hd):(4'ha)]);
            end
          reg517 <= wire75[(4'he):(4'hc)];
          reg518 = (&((reg142[(3'h7):(3'h5)] ?
              reg176[(5'h10):(4'hc)] : $signed(reg86)) + {reg137,
              ($signed(reg186) | reg92)}));
          reg519 <= ($unsigned((~&(&$signed(reg186)))) || (~($unsigned((8'hab)) == reg124)));
        end
      else
        begin
          for (forvar512 = (1'h0); (forvar512 < (1'h0)); forvar512 = (forvar512 + (1'h1)))
            begin
              reg514 <= $signed({($unsigned($unsigned(reg109)) == $unsigned(reg109)),
                  $unsigned(forvar512[(2'h3):(1'h1)])});
              reg516 = $signed((|$unsigned((~|reg137[(1'h1):(1'h1)]))));
              reg517 <= (((reg128[(2'h2):(1'h1)] ?
                          (reg512[(2'h3):(2'h2)] ?
                              $signed(wire76) : reg175[(4'h8):(4'h8)]) : (wire78 << (~reg146))) ?
                      (reg86 && ({(7'h46), reg144} ?
                          (reg144 ?
                              reg123 : (8'hb3)) : (-reg517))) : $unsigned(($signed(reg90) != reg81))) ?
                  ((((reg192 ? reg513 : (8'ha0)) ?
                              (^reg86) : $unsigned(reg92)) ?
                          $unsigned(reg176) : reg512[(5'h10):(3'h7)]) ?
                      {reg188,
                          (~|(~|(8'ha0)))} : reg146[(3'h4):(1'h1)]) : $unsigned(reg175));
              reg518 = ($signed(reg97) ?
                  $signed(reg515) : $signed((~|{$signed(reg180), (+reg511)})));
            end
        end
      reg520 = ((~|reg103[(3'h4):(2'h2)]) ? reg146[(3'h5):(1'h1)] : reg176);
    end
  assign wire521 = $signed((reg177[(2'h3):(1'h0)] ?
                       (reg134[(4'h9):(2'h3)] << (~((8'ha3) ?
                           reg192 : reg122))) : ((~&reg517) <<< $signed($signed((7'h42))))));
  module522 #() modinst655 (wire654, clk, reg90, reg79, reg84, reg142, reg153);
  assign wire656 = $signed(wire77);
  assign wire657 = $unsigned(wire73);
  assign wire658 = reg511;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module522  (y, clk, wire527, wire526, wire525, wire524, wire523);
  output wire [(32'h5f6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire527;
  input wire [(2'h3):(1'h0)] wire526;
  input wire [(5'h12):(1'h0)] wire525;
  input wire [(3'h7):(1'h0)] wire524;
  input wire [(5'h13):(1'h0)] wire523;
  wire signed [(5'h15):(1'h0)] wire651;
  wire signed [(2'h2):(1'h0)] wire650;
  wire [(3'h7):(1'h0)] wire563;
  reg [(3'h7):(1'h0)] reg646 = (1'h0);
  reg [(5'h16):(1'h0)] reg637 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg633 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg632 = (1'h0);
  reg signed [(4'he):(1'h0)] reg631 = (1'h0);
  reg [(4'h9):(1'h0)] reg627 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg626 = (1'h0);
  reg [(4'hb):(1'h0)] reg623 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg622 = (1'h0);
  reg [(4'ha):(1'h0)] reg616 = (1'h0);
  reg [(5'h10):(1'h0)] reg615 = (1'h0);
  reg [(3'h7):(1'h0)] reg613 = (1'h0);
  reg [(2'h2):(1'h0)] reg611 = (1'h0);
  reg [(4'hb):(1'h0)] reg610 = (1'h0);
  reg [(4'hb):(1'h0)] reg606 = (1'h0);
  reg [(4'ha):(1'h0)] reg601 = (1'h0);
  reg [(3'h4):(1'h0)] reg597 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg592 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg589 = (1'h0);
  reg [(2'h3):(1'h0)] reg587 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg584 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg581 = (1'h0);
  reg [(3'h4):(1'h0)] reg579 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg578 = (1'h0);
  reg [(2'h2):(1'h0)] reg575 = (1'h0);
  reg [(5'h12):(1'h0)] reg574 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg573 = (1'h0);
  reg [(3'h5):(1'h0)] reg571 = (1'h0);
  reg [(5'h10):(1'h0)] reg567 = (1'h0);
  reg signed [(4'he):(1'h0)] reg566 = (1'h0);
  reg [(3'h4):(1'h0)] reg562 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg559 = (1'h0);
  reg [(5'h10):(1'h0)] reg558 = (1'h0);
  reg [(5'h13):(1'h0)] reg554 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg548 = (1'h0);
  reg [(3'h4):(1'h0)] reg541 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg536 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg530 = (1'h0);
  reg [(2'h3):(1'h0)] reg533 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg531 = (1'h0);
  reg [(5'h16):(1'h0)] reg528 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg653 = (1'h0);
  reg [(5'h16):(1'h0)] reg652 = (1'h0);
  reg [(4'ha):(1'h0)] reg649 = (1'h0);
  reg [(5'h12):(1'h0)] forvar641 = (1'h0);
  reg [(3'h6):(1'h0)] reg648 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg647 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg645 = (1'h0);
  reg [(5'h18):(1'h0)] reg644 = (1'h0);
  reg [(4'he):(1'h0)] reg643 = (1'h0);
  reg [(3'h6):(1'h0)] reg642 = (1'h0);
  reg [(2'h3):(1'h0)] reg641 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg640 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar639 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg638 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar636 = (1'h0);
  reg [(5'h12):(1'h0)] reg635 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg634 = (1'h0);
  reg [(5'h11):(1'h0)] reg630 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar629 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg628 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar625 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg624 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar621 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg620 = (1'h0);
  reg [(5'h16):(1'h0)] reg619 = (1'h0);
  reg [(4'hf):(1'h0)] reg618 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg617 = (1'h0);
  reg [(4'ha):(1'h0)] forvar614 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg612 = (1'h0);
  reg [(5'h11):(1'h0)] reg609 = (1'h0);
  reg [(5'h10):(1'h0)] reg608 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg607 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg605 = (1'h0);
  reg [(4'he):(1'h0)] reg604 = (1'h0);
  reg [(4'h9):(1'h0)] reg603 = (1'h0);
  reg [(4'ha):(1'h0)] reg602 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg599 = (1'h0);
  reg [(4'hc):(1'h0)] reg598 = (1'h0);
  reg [(4'hf):(1'h0)] forvar593 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg596 = (1'h0);
  reg [(4'hb):(1'h0)] reg595 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg594 = (1'h0);
  reg [(4'h9):(1'h0)] reg593 = (1'h0);
  reg [(3'h5):(1'h0)] reg591 = (1'h0);
  reg [(3'h7):(1'h0)] reg590 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg588 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar586 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg585 = (1'h0);
  reg [(4'h9):(1'h0)] forvar583 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg582 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg580 = (1'h0);
  reg [(5'h11):(1'h0)] forvar577 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg576 = (1'h0);
  reg [(2'h3):(1'h0)] reg572 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg570 = (1'h0);
  reg [(4'ha):(1'h0)] reg569 = (1'h0);
  reg [(4'hd):(1'h0)] reg568 = (1'h0);
  reg [(5'h15):(1'h0)] reg565 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar564 = (1'h0);
  reg [(3'h7):(1'h0)] forvar561 = (1'h0);
  reg [(5'h11):(1'h0)] reg560 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar557 = (1'h0);
  reg [(4'ha):(1'h0)] reg556 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg555 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg553 = (1'h0);
  reg [(3'h6):(1'h0)] reg552 = (1'h0);
  reg [(4'hd):(1'h0)] forvar551 = (1'h0);
  reg [(2'h2):(1'h0)] reg550 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg549 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg547 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar546 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg545 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar544 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg543 = (1'h0);
  reg [(4'hf):(1'h0)] reg542 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg540 = (1'h0);
  reg [(5'h15):(1'h0)] reg539 = (1'h0);
  reg [(4'ha):(1'h0)] forvar538 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg537 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg534 = (1'h0);
  reg [(4'h8):(1'h0)] reg532 = (1'h0);
  reg [(3'h7):(1'h0)] forvar530 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg529 = (1'h0);
  assign y = {wire651,
                 wire650,
                 wire563,
                 reg646,
                 reg637,
                 reg633,
                 reg632,
                 reg631,
                 reg627,
                 reg626,
                 reg623,
                 reg622,
                 reg616,
                 reg615,
                 reg613,
                 reg611,
                 reg610,
                 reg606,
                 reg601,
                 reg597,
                 reg592,
                 reg589,
                 reg587,
                 reg584,
                 reg581,
                 reg579,
                 reg578,
                 reg575,
                 reg574,
                 reg573,
                 reg571,
                 reg567,
                 reg566,
                 reg562,
                 reg559,
                 reg558,
                 reg554,
                 reg548,
                 reg541,
                 reg536,
                 reg530,
                 reg533,
                 reg531,
                 reg528,
                 reg653,
                 reg652,
                 reg649,
                 forvar641,
                 reg648,
                 reg647,
                 reg645,
                 reg644,
                 reg643,
                 reg642,
                 reg641,
                 reg640,
                 forvar639,
                 reg638,
                 forvar636,
                 reg635,
                 reg634,
                 reg630,
                 forvar629,
                 reg628,
                 forvar625,
                 reg624,
                 forvar621,
                 reg620,
                 reg619,
                 reg618,
                 reg617,
                 forvar614,
                 reg612,
                 reg609,
                 reg608,
                 reg607,
                 reg605,
                 reg604,
                 reg603,
                 reg602,
                 reg600,
                 reg599,
                 reg598,
                 forvar593,
                 reg596,
                 reg595,
                 reg594,
                 reg593,
                 reg591,
                 reg590,
                 reg588,
                 forvar586,
                 reg585,
                 forvar583,
                 reg582,
                 reg580,
                 forvar577,
                 reg576,
                 reg572,
                 reg570,
                 reg569,
                 reg568,
                 reg565,
                 forvar564,
                 forvar561,
                 reg560,
                 forvar557,
                 reg556,
                 reg555,
                 reg553,
                 reg552,
                 forvar551,
                 reg550,
                 reg549,
                 reg547,
                 forvar546,
                 reg545,
                 forvar544,
                 reg543,
                 reg542,
                 reg540,
                 reg539,
                 forvar538,
                 reg537,
                 reg535,
                 reg534,
                 reg532,
                 forvar530,
                 reg529,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire525[(3'h5):(1'h0)])
        begin
          reg528 <= {(($unsigned((wire525 ? (8'had) : (7'h48))) ?
                  wire525 : ((wire524 ?
                      wire526 : wire527) & {wire524})) >>> $unsigned(({wire525,
                      wire526} ?
                  (wire527 << (8'h9d)) : (wire527 + wire523)))),
              wire526[(1'h0):(1'h0)]};
          reg529 = wire526[(1'h0):(1'h0)];
          for (forvar530 = (1'h0); (forvar530 < (2'h2)); forvar530 = (forvar530 + (1'h1)))
            begin
              reg531 <= ($signed(($unsigned(forvar530[(1'h1):(1'h1)]) ?
                  ({reg529} ? {wire525, reg529} : (|wire527)) : (~^(wire527 ?
                      wire525 : wire524)))) != (^~({$unsigned((8'hbf)),
                      $signed(wire525)} ?
                  wire523[(1'h0):(1'h0)] : $signed(wire527[(2'h2):(2'h2)]))));
              reg532 = $unsigned(wire523[(4'hc):(4'hb)]);
              reg533 <= reg532[(1'h0):(1'h0)];
              reg534 = ($unsigned((^(-(reg531 ? reg533 : (8'hb4))))) ?
                  (wire525 ^ ($unsigned(reg529) ?
                      ((forvar530 ? reg533 : wire527) ?
                          $signed((8'ha7)) : reg533[(2'h3):(2'h2)]) : wire524[(1'h1):(1'h0)])) : reg532);
            end
          reg535 = forvar530;
        end
      else
        begin
          if ((((8'hbb) << ($signed(forvar530) ?
              ($signed((8'ha1)) ?
                  (!wire524) : ((8'hb1) >>> reg529)) : reg529)) * $signed(wire527)))
            begin
              reg529 = (8'ha6);
              reg530 <= $unsigned($unsigned(((reg534 ?
                      $unsigned(reg528) : (8'hb5)) ?
                  (wire527 < (+wire527)) : reg533)));
              reg532 = (-$unsigned($unsigned($signed(reg532[(2'h3):(2'h2)]))));
              reg534 = (~^reg532[(2'h2):(2'h2)]);
              reg535 = wire524[(3'h7):(3'h6)];
            end
          else
            begin
              reg528 <= reg529[(3'h4):(2'h3)];
            end
          reg536 <= (((~^($unsigned(wire527) >= (reg534 ?
              wire526 : (8'hab)))) >= wire527) ^ $signed(($unsigned(reg528) <<< $signed((8'hb1)))));
          reg537 = ((+$unsigned(((wire525 != (8'ha4)) - $unsigned(reg531)))) - $unsigned(((reg535 + (reg532 <<< (8'hbb))) < ($unsigned(reg531) ?
              (reg529 ? reg532 : reg529) : ((8'ha5) ? reg534 : (8'h9e))))));
          for (forvar538 = (1'h0); (forvar538 < (1'h1)); forvar538 = (forvar538 + (1'h1)))
            begin
              reg539 = reg528;
              reg540 = (+($signed((forvar538[(2'h3):(1'h0)] ?
                      wire524[(3'h4):(2'h3)] : (^~reg535))) ?
                  forvar538 : ($signed({reg534}) ?
                      wire523[(4'hc):(4'hb)] : ($unsigned(wire523) ?
                          reg536[(3'h5):(2'h3)] : wire526[(2'h2):(2'h2)]))));
              reg541 <= reg531;
              reg542 = (wire527 <<< reg532);
            end
          reg543 = reg532[(3'h7):(3'h6)];
        end
      for (forvar544 = (1'h0); (forvar544 < (3'h4)); forvar544 = (forvar544 + (1'h1)))
        begin
          reg545 = ($unsigned(forvar538) ?
              $unsigned(reg531) : {{{(reg537 ? (8'h9d) : reg532)},
                      ($signed(reg530) ? $signed(reg532) : reg540)}});
          for (forvar546 = (1'h0); (forvar546 < (2'h3)); forvar546 = (forvar546 + (1'h1)))
            begin
              reg547 = ((((~|reg537[(3'h6):(3'h5)]) ~^ ((reg535 & reg539) ?
                  (reg541 ~^ reg532) : reg528[(3'h7):(3'h6)])) | $unsigned({wire524,
                  $signed(reg532)})) <<< $signed(((-((7'h49) << reg539)) ?
                  ({forvar530} ? $signed((7'h40)) : (~&reg539)) : reg536)));
              reg548 <= $signed($signed($signed(forvar530[(3'h6):(3'h5)])));
              reg549 = (((reg548 <<< $unsigned($unsigned(wire524))) * (reg536[(4'h8):(2'h2)] ?
                      reg547[(1'h0):(1'h0)] : ($signed(forvar546) <<< (reg532 < reg543)))) ?
                  (-reg537) : wire527);
              reg550 = $signed($signed((~^(&$signed(wire526)))));
            end
          for (forvar551 = (1'h0); (forvar551 < (1'h0)); forvar551 = (forvar551 + (1'h1)))
            begin
              reg552 = {reg549[(4'hd):(4'hc)], reg543[(4'h8):(3'h6)]};
              reg553 = reg543[(1'h0):(1'h0)];
              reg554 <= ((wire526 ?
                      (forvar551 <= ({reg545} == (reg553 ?
                          reg539 : (8'h9e)))) : (~&reg545)) ?
                  (~($unsigned(forvar538) > (~|(wire524 ?
                      (8'ha6) : reg547)))) : $unsigned(reg537[(3'h6):(1'h1)]));
              reg555 = (({(^reg548[(2'h3):(1'h1)]),
                  $unsigned((reg529 <<< wire527))} == (^(^(reg535 ?
                  reg542 : reg540)))) || reg543[(2'h3):(2'h3)]);
            end
          reg556 = {$signed($unsigned(forvar538[(4'ha):(4'h8)]))};
          for (forvar557 = (1'h0); (forvar557 < (2'h3)); forvar557 = (forvar557 + (1'h1)))
            begin
              reg558 <= $signed((((&(8'hb8)) ?
                  ((reg555 ? reg555 : reg555) ?
                      (^reg552) : (wire525 ? wire524 : (8'ha7))) : ((reg530 ?
                      reg545 : reg542) ^~ $signed(reg543))) ~^ $unsigned((~&$unsigned(wire525)))));
              reg559 <= $unsigned({(reg558[(4'h8):(1'h1)] ~^ $signed({reg537})),
                  reg541});
              reg560 = (($unsigned((-(reg548 ?
                  forvar546 : (8'h9d)))) > (reg547[(4'h9):(1'h0)] ^~ ($signed(reg542) ?
                  {reg536} : (reg549 ? reg554 : (8'ha6))))) << (~(reg554 ?
                  reg531 : (|(reg543 * forvar551)))));
            end
        end
      for (forvar561 = (1'h0); (forvar561 < (3'h4)); forvar561 = (forvar561 + (1'h1)))
        begin
          reg562 <= ((|(((^~reg545) || $signed(reg556)) ? {reg530} : reg553)) ?
              reg534[(4'h8):(3'h6)] : (~|reg532[(1'h1):(1'h0)]));
        end
    end
  assign wire563 = reg558[(3'h7):(1'h1)];
  always
    @(posedge clk) begin
      for (forvar564 = (1'h0); (forvar564 < (1'h1)); forvar564 = (forvar564 + (1'h1)))
        begin
          reg565 = reg528;
          reg566 <= $unsigned($unsigned((~&$unsigned(reg533[(2'h3):(1'h1)]))));
          reg567 <= forvar564[(2'h3):(2'h3)];
          reg568 = ((reg528[(5'h13):(2'h2)] ?
              $unsigned($signed(((8'hbc) <= (8'h9e)))) : $signed(reg533)) >= (|$signed(reg536[(4'he):(4'hb)])));
          if (reg528[(5'h13):(3'h7)])
            begin
              reg569 = $unsigned($unsigned($unsigned($unsigned({reg568,
                  wire524}))));
              reg570 = $unsigned(($unsigned($unsigned(reg533[(1'h0):(1'h0)])) <<< $unsigned(reg559)));
              reg571 <= {$unsigned($signed(wire523[(4'hf):(4'h8)])),
                  (($signed($signed(wire525)) > $unsigned({reg548})) ^~ reg533[(1'h0):(1'h0)])};
              reg572 = (|wire525);
              reg573 <= ($signed(wire525) >= ($unsigned(reg541[(2'h3):(1'h0)]) | reg569));
            end
          else
            begin
              reg569 = wire523;
              reg570 = {$unsigned(reg566[(4'hc):(4'h8)]), reg573};
              reg571 <= (+((~^(~|reg562)) ?
                  reg530 : $signed($unsigned({reg571}))));
              reg572 = $unsigned((reg536[(1'h1):(1'h0)] || wire526[(1'h0):(1'h0)]));
            end
        end
      reg574 <= {((~&(&$unsigned(forvar564))) ?
              reg571[(2'h3):(1'h0)] : (reg530 ?
                  $signed((~^reg567)) : ($unsigned(reg568) <= wire563))),
          reg533[(2'h3):(2'h2)]};
      if ((~$signed({wire527, $unsigned($unsigned(reg554))})))
        begin
          reg575 <= ($unsigned((({wire526, reg570} ?
                  (~reg530) : reg573) << (8'haa))) ?
              reg569[(1'h0):(1'h0)] : $unsigned(reg571));
          reg576 = (reg531 * reg559[(1'h1):(1'h1)]);
        end
      else
        begin
          reg576 = ($signed((+reg571[(1'h0):(1'h0)])) >> ($signed($signed($signed(wire523))) * (7'h48)));
          for (forvar577 = (1'h0); (forvar577 < (1'h1)); forvar577 = (forvar577 + (1'h1)))
            begin
              reg578 <= $unsigned({(|reg559[(1'h0):(1'h0)]),
                  $unsigned(({wire527, reg558} ?
                      ((7'h45) | reg559) : reg559[(3'h6):(1'h0)]))});
              reg579 <= reg568;
              reg580 = (wire523 ?
                  (^reg570[(2'h3):(1'h1)]) : $signed({($signed(wire563) <<< reg579[(1'h0):(1'h0)]),
                      (7'h42)}));
              reg581 <= (7'h46);
              reg582 = ({(($signed(reg531) > (reg565 ?
                      reg558 : reg575)) ~^ ((reg571 ? reg565 : (8'hb1)) ?
                      wire526[(2'h3):(1'h0)] : $unsigned(reg570)))} || $signed($signed(reg581[(1'h0):(1'h0)])));
            end
          for (forvar583 = (1'h0); (forvar583 < (1'h0)); forvar583 = (forvar583 + (1'h1)))
            begin
              reg584 <= ({(&({(8'hb3)} ?
                          reg573[(2'h3):(1'h0)] : (reg558 - reg568)))} ?
                  (|$unsigned({reg554[(4'hc):(4'hb)],
                      (reg559 == reg531)})) : reg579[(1'h0):(1'h0)]);
            end
        end
      reg585 = (reg533 ?
          reg531 : (($signed((reg576 ? wire523 : wire525)) ?
              $unsigned($unsigned(reg531)) : (^reg554)) >>> $signed((+(8'haf)))));
      if ((~|((8'hb5) ? reg567 : (+$unsigned((reg566 <<< wire527))))))
        begin
          for (forvar586 = (1'h0); (forvar586 < (2'h3)); forvar586 = (forvar586 + (1'h1)))
            begin
              reg587 <= $unsigned(reg559);
              reg588 = $unsigned($signed(reg568[(1'h1):(1'h0)]));
              reg589 <= ((($signed((~&reg562)) || ($unsigned(reg578) && ((8'hbc) >>> (8'h9c)))) != ($signed(reg578[(1'h0):(1'h0)]) > $unsigned(reg558[(4'h9):(3'h7)]))) ?
                  $unsigned((^(8'hbc))) : (~&$signed($unsigned($unsigned(forvar583)))));
            end
          if ({$unsigned($unsigned($unsigned(((7'h47) <<< reg554)))),
              $signed(wire525[(4'h9):(3'h4)])})
            begin
              reg590 = $unsigned(wire525[(2'h2):(1'h1)]);
              reg591 = reg574;
              reg592 <= wire563;
            end
          else
            begin
              reg590 = wire527;
              reg591 = (^((reg573 ?
                      $signed((reg541 ?
                          reg579 : reg566)) : ((~^reg536) && wire523)) ?
                  reg585 : $unsigned($unsigned($unsigned(reg566)))));
              reg593 = ((&(reg589[(2'h3):(1'h0)] ?
                  (((8'ha9) < reg575) ~^ $unsigned(reg536)) : ((reg579 ?
                          reg573 : wire527) ?
                      wire525 : (forvar577 - reg566)))) <= reg568);
              reg594 = reg530[(3'h5):(3'h4)];
              reg595 = $unsigned(reg567[(4'hf):(3'h6)]);
            end
          reg596 = ($signed(reg569) ? reg587 : reg592[(3'h4):(3'h4)]);
          reg597 <= (reg590 > ((8'ha3) ?
              ($unsigned(reg562) >= $unsigned($unsigned(reg589))) : reg533));
        end
      else
        begin
          for (forvar586 = (1'h0); (forvar586 < (1'h0)); forvar586 = (forvar586 + (1'h1)))
            begin
              reg588 = {reg597, reg566[(3'h7):(1'h0)]};
              reg589 <= reg559;
              reg592 <= reg541;
            end
          for (forvar593 = (1'h0); (forvar593 < (1'h0)); forvar593 = (forvar593 + (1'h1)))
            begin
              reg597 <= reg567[(4'h9):(1'h0)];
              reg598 = {(((reg541[(1'h0):(1'h0)] ?
                              $unsigned(wire527) : (reg570 ?
                                  forvar564 : reg531)) ?
                          ((!forvar593) || (reg579 ?
                              (7'h42) : reg579)) : ($unsigned((8'hbd)) & $unsigned(reg530))) ?
                      reg584 : $unsigned((wire524 ^~ wire563[(3'h5):(3'h4)]))),
                  (~{((~&reg579) ?
                          forvar564[(3'h4):(1'h0)] : $signed(forvar586))})};
              reg599 = reg574;
            end
          reg600 = $signed({(-(8'ha9)), $signed(($signed(reg572) && (8'hb0)))});
        end
    end
  always
    @(posedge clk) begin
      reg601 <= $signed((-reg581));
      if ($unsigned(reg558))
        begin
          reg602 = $unsigned($signed(($signed(reg531) ?
              $unsigned((&reg528)) : wire524)));
          if ({$signed(reg558[(3'h4):(1'h1)]), reg579})
            begin
              reg603 = reg562[(2'h2):(1'h0)];
              reg604 = (~&(~reg592));
              reg605 = reg533;
            end
          else
            begin
              reg606 <= {({$unsigned((reg548 ? wire523 : reg584)),
                          ($signed(reg530) ? {wire524} : {reg536, reg581})} ?
                      {reg574} : {(reg604 ?
                              ((8'h9c) <<< wire524) : (-reg574))}),
                  reg581[(2'h3):(2'h3)]};
              reg607 = (reg581[(3'h7):(1'h0)] ?
                  (reg575 ?
                      {(reg528[(3'h4):(2'h3)] ?
                              reg567 : (reg587 < reg562))} : reg602[(4'ha):(4'ha)]) : (-(|$unsigned($unsigned(reg602)))));
              reg608 = (~&{(reg554[(5'h10):(4'hd)] + ({(8'ha8), (8'hbc)} ?
                      $unsigned(reg574) : reg530)),
                  reg554[(5'h12):(1'h0)]});
              reg609 = $unsigned(wire563[(3'h4):(3'h4)]);
            end
          reg610 <= (reg609 ?
              ((((reg604 ? reg536 : reg607) ?
                  $unsigned(wire563) : reg578) >> ((reg604 ? reg587 : reg603) ?
                  (wire563 ? reg573 : wire523) : reg528)) << {(reg530 ?
                      (|(8'hac)) : reg574),
                  $signed(reg541[(2'h3):(1'h1)])}) : $unsigned($unsigned(wire563)));
          reg611 <= (reg571 < reg578[(4'hf):(3'h4)]);
        end
      else
        begin
          if ((~^$unsigned((reg567 ?
              (^(wire524 ? reg605 : wire523)) : reg587[(1'h1):(1'h1)]))))
            begin
              reg602 = ((!(wire563[(2'h2):(1'h1)] ?
                  reg536[(5'h10):(1'h0)] : $signed(reg562))) ~^ (~|($unsigned((^reg566)) ?
                  reg573 : reg605[(5'h14):(5'h14)])));
            end
          else
            begin
              reg606 <= reg584[(5'h10):(4'hc)];
              reg607 = $signed($signed((((~^reg604) | (~&reg575)) ?
                  ((reg528 >>> reg567) < reg606[(3'h5):(2'h3)]) : ((^~reg609) ?
                      (reg530 ~^ reg573) : reg574[(3'h6):(3'h6)]))));
              reg610 <= (((~reg597[(2'h2):(1'h0)]) ^ {(reg554[(4'h9):(4'h8)] ~^ $signed(wire526)),
                      ((reg589 ^ reg604) - $signed((8'hbe)))}) ?
                  reg554[(5'h10):(4'h9)] : (reg605[(4'ha):(4'h9)] ?
                      ($signed($signed(reg571)) ?
                          (!(8'hb7)) : $signed(wire527)) : $signed(($unsigned((8'hb8)) ~^ reg607[(4'ha):(3'h5)]))));
            end
        end
      reg612 = (^~(8'hae));
      reg613 <= $unsigned((8'h9d));
    end
  always
    @(posedge clk) begin
      for (forvar614 = (1'h0); (forvar614 < (2'h3)); forvar614 = (forvar614 + (1'h1)))
        begin
          if ($unsigned(reg559))
            begin
              reg615 <= $unsigned($signed(reg574[(4'h8):(3'h5)]));
              reg616 <= $signed(((((^~reg592) ?
                  $unsigned(wire525) : (reg613 ~^ reg592)) > (!reg597)) && $signed((!{reg548,
                  reg589}))));
              reg617 = reg573[(1'h0):(1'h0)];
              reg618 = reg558[(4'hc):(1'h1)];
            end
          else
            begin
              reg615 <= (+(~&(!reg579)));
              reg617 = (($unsigned($signed($unsigned(reg617))) || (($signed((7'h46)) ^ (8'hab)) << ($unsigned(reg617) & (reg581 ?
                      reg597 : reg530)))) ?
                  reg559[(1'h0):(1'h0)] : ({{wire526[(1'h0):(1'h0)],
                              (reg559 ? reg601 : (8'hb2))}} ?
                      (wire525[(3'h5):(2'h3)] ?
                          $signed($signed((8'hba))) : ($unsigned(reg531) - $unsigned((7'h40)))) : reg578[(2'h3):(2'h2)]));
              reg618 = $unsigned((reg530[(5'h10):(4'hb)] ^ (reg566[(4'ha):(4'ha)] & (^reg613))));
              reg619 = $unsigned(((^~($unsigned(reg567) + $signed((8'hbd)))) ~^ reg581));
              reg620 = (8'ha9);
            end
          for (forvar621 = (1'h0); (forvar621 < (2'h3)); forvar621 = (forvar621 + (1'h1)))
            begin
              reg622 <= (+(reg530 ? wire563 : (reg619 ? {reg615} : reg589)));
              reg623 <= (($signed(reg536[(4'ha):(1'h1)]) ^~ {(!(^(8'hbc))),
                  wire523[(4'h9):(3'h4)]}) || ({$unsigned({reg536,
                      reg617})} != (!reg587[(2'h3):(2'h2)])));
              reg624 = ((reg597 ?
                  (|(&{reg530})) : reg574[(5'h10):(1'h1)]) || (~|(reg530 & $signed(reg541[(1'h1):(1'h0)]))));
            end
          for (forvar625 = (1'h0); (forvar625 < (3'h4)); forvar625 = (forvar625 + (1'h1)))
            begin
              reg626 <= (reg559 << $signed($signed(reg618[(4'hd):(2'h2)])));
              reg627 <= wire525[(3'h5):(2'h3)];
              reg628 = $unsigned($signed($unsigned($signed(reg623[(1'h1):(1'h1)]))));
            end
          for (forvar629 = (1'h0); (forvar629 < (1'h0)); forvar629 = (forvar629 + (1'h1)))
            begin
              reg630 = {{($unsigned(reg622) ?
                          wire524[(1'h1):(1'h0)] : (^{reg615, reg558}))}};
              reg631 <= $signed((~&reg592));
              reg632 <= (~^{reg548});
            end
        end
      reg633 <= {$unsigned(reg533)};
      reg634 = reg610;
      reg635 = (8'ha2);
      for (forvar636 = (1'h0); (forvar636 < (1'h1)); forvar636 = (forvar636 + (1'h1)))
        begin
          reg637 <= $signed(((($signed(reg562) > $signed(reg573)) & $unsigned((forvar625 ?
                  reg613 : forvar629))) ?
              ({$signed(reg548), (forvar629 && wire527)} ?
                  $signed((&reg541)) : (8'hb2)) : $signed((^(^reg558)))));
        end
    end
  always
    @(posedge clk) begin
      reg638 = reg633[(2'h2):(1'h1)];
      for (forvar639 = (1'h0); (forvar639 < (1'h0)); forvar639 = (forvar639 + (1'h1)))
        begin
          reg640 = (+reg533);
        end
      if ($signed(reg530))
        begin
          reg641 = $unsigned(reg578);
          if ($unsigned((((reg638 <= wire523) ?
                  (8'hbc) : $signed(reg641[(1'h0):(1'h0)])) ?
              (((reg587 ? reg571 : reg562) == (&reg533)) ?
                  reg579[(3'h4):(2'h3)] : ((-reg623) ?
                      reg571 : (reg611 && reg592))) : wire523)))
            begin
              reg642 = (reg559[(2'h3):(2'h3)] ^ ((8'hac) ?
                  reg530 : (reg592[(3'h6):(1'h1)] == ((reg558 && (8'ha9)) >>> reg531[(1'h1):(1'h1)]))));
              reg643 = reg578;
              reg644 = $unsigned(reg574[(4'hf):(4'he)]);
              reg645 = ((|$unsigned($signed($unsigned((8'ha7))))) ?
                  wire563 : (reg548 ?
                      (8'ha6) : (wire526[(2'h3):(1'h0)] ?
                          $unsigned(reg589) : ({reg530, (8'ha6)} ?
                              {reg567, reg567} : reg640))));
            end
          else
            begin
              reg646 <= (($signed({$unsigned(reg575)}) << $signed($unsigned((reg641 ?
                  reg645 : reg566)))) >> (|reg637));
              reg647 = {(!reg642[(1'h0):(1'h0)]),
                  (($signed(reg643) << ($signed(forvar639) >= (7'h40))) >> {{(reg548 ~^ reg554),
                          reg554[(2'h2):(2'h2)]},
                      ((reg554 ? (8'hb7) : reg597) ?
                          $signed(reg640) : (reg616 < (8'hb1)))})};
            end
          reg648 = wire526;
        end
      else
        begin
          for (forvar641 = (1'h0); (forvar641 < (2'h3)); forvar641 = (forvar641 + (1'h1)))
            begin
              reg642 = (~^$unsigned($unsigned($unsigned($signed(reg643)))));
            end
        end
      reg649 = $unsigned(reg533);
    end
  assign wire650 = (~(reg574[(5'h11):(1'h1)] ?
                       (reg615[(2'h3):(2'h2)] ?
                           $unsigned(reg592) : (^~wire526[(1'h0):(1'h0)])) : $signed((^reg530[(1'h0):(1'h0)]))));
  assign wire651 = ((reg548 + (!$unsigned($unsigned(reg528)))) >> $signed(wire526));
  always
    @(posedge clk) begin
      reg652 = {(~|({(&wire524)} ^~ $signed($unsigned((7'h49)))))};
      reg653 = (8'h9f);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module195  (y, clk, wire199, wire198, wire197, wire196);
  output wire [(32'h1093):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire199;
  input wire [(4'hc):(1'h0)] wire198;
  input wire signed [(5'h15):(1'h0)] wire197;
  input wire signed [(5'h12):(1'h0)] wire196;
  wire [(4'hf):(1'h0)] wire507;
  wire signed [(4'h8):(1'h0)] wire424;
  wire [(4'hb):(1'h0)] wire324;
  wire signed [(5'h15):(1'h0)] wire249;
  wire signed [(5'h11):(1'h0)] wire248;
  wire [(5'h15):(1'h0)] wire247;
  wire signed [(5'h16):(1'h0)] wire226;
  wire signed [(4'hc):(1'h0)] wire225;
  wire signed [(4'ha):(1'h0)] wire224;
  reg signed [(5'h12):(1'h0)] reg490 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg504 = (1'h0);
  reg [(2'h2):(1'h0)] reg502 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg501 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg496 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg495 = (1'h0);
  reg [(5'h14):(1'h0)] reg493 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg488 = (1'h0);
  reg [(2'h3):(1'h0)] reg485 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg482 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg481 = (1'h0);
  reg [(4'ha):(1'h0)] reg480 = (1'h0);
  reg [(5'h17):(1'h0)] reg476 = (1'h0);
  reg [(4'hc):(1'h0)] reg473 = (1'h0);
  reg [(3'h5):(1'h0)] reg472 = (1'h0);
  reg [(4'he):(1'h0)] reg471 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg470 = (1'h0);
  reg [(4'h9):(1'h0)] reg469 = (1'h0);
  reg [(3'h6):(1'h0)] reg466 = (1'h0);
  reg [(4'hb):(1'h0)] reg460 = (1'h0);
  reg [(2'h2):(1'h0)] reg457 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg456 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg455 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg453 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg451 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg450 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg449 = (1'h0);
  reg [(5'h10):(1'h0)] reg447 = (1'h0);
  reg [(5'h18):(1'h0)] reg446 = (1'h0);
  reg [(4'he):(1'h0)] reg441 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg440 = (1'h0);
  reg [(2'h3):(1'h0)] reg438 = (1'h0);
  reg [(2'h2):(1'h0)] reg436 = (1'h0);
  reg [(3'h6):(1'h0)] reg435 = (1'h0);
  reg [(2'h3):(1'h0)] reg434 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg432 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg430 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg428 = (1'h0);
  reg [(4'ha):(1'h0)] reg427 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg426 = (1'h0);
  reg signed [(4'he):(1'h0)] reg423 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg422 = (1'h0);
  reg [(5'h15):(1'h0)] reg421 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg418 = (1'h0);
  reg [(4'hc):(1'h0)] reg415 = (1'h0);
  reg [(4'hf):(1'h0)] reg413 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg409 = (1'h0);
  reg [(3'h5):(1'h0)] reg408 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg405 = (1'h0);
  reg [(5'h15):(1'h0)] reg404 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg401 = (1'h0);
  reg [(5'h10):(1'h0)] reg400 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg399 = (1'h0);
  reg [(5'h14):(1'h0)] reg398 = (1'h0);
  reg [(4'he):(1'h0)] reg397 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg396 = (1'h0);
  reg [(4'hb):(1'h0)] reg392 = (1'h0);
  reg [(3'h7):(1'h0)] reg390 = (1'h0);
  reg [(4'hf):(1'h0)] reg388 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg376 = (1'h0);
  reg [(4'hb):(1'h0)] reg373 = (1'h0);
  reg [(5'h13):(1'h0)] reg372 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg371 = (1'h0);
  reg [(4'hf):(1'h0)] reg370 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg366 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg365 = (1'h0);
  reg [(4'h8):(1'h0)] reg364 = (1'h0);
  reg [(4'h9):(1'h0)] reg363 = (1'h0);
  reg [(5'h15):(1'h0)] reg362 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg360 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg353 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg352 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg351 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg349 = (1'h0);
  reg [(3'h7):(1'h0)] reg346 = (1'h0);
  reg [(4'hb):(1'h0)] reg345 = (1'h0);
  reg [(4'hb):(1'h0)] reg343 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg342 = (1'h0);
  reg [(2'h2):(1'h0)] reg339 = (1'h0);
  reg [(4'h8):(1'h0)] reg338 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg333 = (1'h0);
  reg [(5'h14):(1'h0)] reg336 = (1'h0);
  reg [(5'h10):(1'h0)] reg334 = (1'h0);
  reg [(5'h12):(1'h0)] reg329 = (1'h0);
  reg [(5'h17):(1'h0)] reg326 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg313 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg323 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg322 = (1'h0);
  reg [(5'h10):(1'h0)] reg320 = (1'h0);
  reg [(5'h10):(1'h0)] reg316 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg310 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg307 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg306 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg304 = (1'h0);
  reg [(3'h4):(1'h0)] reg303 = (1'h0);
  reg [(4'he):(1'h0)] reg302 = (1'h0);
  reg [(2'h2):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg299 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg298 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg297 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg284 = (1'h0);
  reg [(5'h13):(1'h0)] reg282 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg280 = (1'h0);
  reg [(4'h9):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg275 = (1'h0);
  reg [(4'h9):(1'h0)] reg273 = (1'h0);
  reg [(4'hb):(1'h0)] reg270 = (1'h0);
  reg [(5'h12):(1'h0)] reg267 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg266 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg263 = (1'h0);
  reg [(5'h15):(1'h0)] reg262 = (1'h0);
  reg [(5'h13):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg257 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg256 = (1'h0);
  reg [(4'hb):(1'h0)] reg254 = (1'h0);
  reg [(5'h14):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg244 = (1'h0);
  reg [(4'he):(1'h0)] reg242 = (1'h0);
  reg [(4'hf):(1'h0)] reg238 = (1'h0);
  reg [(5'h16):(1'h0)] reg237 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg234 = (1'h0);
  reg [(4'hb):(1'h0)] reg231 = (1'h0);
  reg [(5'h16):(1'h0)] reg230 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg227 = (1'h0);
  reg [(4'h9):(1'h0)] reg223 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg214 = (1'h0);
  reg [(5'h12):(1'h0)] reg210 = (1'h0);
  reg [(5'h18):(1'h0)] reg204 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg203 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg202 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg201 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg497 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar496 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg494 = (1'h0);
  reg [(4'hb):(1'h0)] forvar491 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg506 = (1'h0);
  reg [(4'hf):(1'h0)] reg505 = (1'h0);
  reg [(3'h4):(1'h0)] forvar503 = (1'h0);
  reg [(4'ha):(1'h0)] reg500 = (1'h0);
  reg [(4'ha):(1'h0)] reg499 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg498 = (1'h0);
  reg [(5'h10):(1'h0)] forvar497 = (1'h0);
  reg [(4'h8):(1'h0)] forvar494 = (1'h0);
  reg [(3'h6):(1'h0)] reg492 = (1'h0);
  reg [(5'h17):(1'h0)] reg491 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar490 = (1'h0);
  reg [(4'hd):(1'h0)] reg489 = (1'h0);
  reg [(3'h7):(1'h0)] reg487 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg486 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg484 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg483 = (1'h0);
  reg [(5'h15):(1'h0)] reg479 = (1'h0);
  reg signed [(4'he):(1'h0)] reg478 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar477 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg475 = (1'h0);
  reg [(5'h16):(1'h0)] reg474 = (1'h0);
  reg [(5'h13):(1'h0)] reg468 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg467 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg465 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar452 = (1'h0);
  reg [(5'h16):(1'h0)] reg464 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg463 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg462 = (1'h0);
  reg [(3'h7):(1'h0)] reg461 = (1'h0);
  reg [(4'hb):(1'h0)] reg459 = (1'h0);
  reg [(4'h9):(1'h0)] forvar458 = (1'h0);
  reg [(4'hf):(1'h0)] reg454 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg452 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg448 = (1'h0);
  reg [(5'h18):(1'h0)] forvar445 = (1'h0);
  reg [(3'h5):(1'h0)] reg444 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar443 = (1'h0);
  reg [(4'hb):(1'h0)] forvar442 = (1'h0);
  reg [(5'h14):(1'h0)] forvar434 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar425 = (1'h0);
  reg [(5'h16):(1'h0)] reg439 = (1'h0);
  reg [(4'he):(1'h0)] reg437 = (1'h0);
  reg [(4'he):(1'h0)] reg433 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg431 = (1'h0);
  reg [(5'h18):(1'h0)] reg429 = (1'h0);
  reg [(3'h5):(1'h0)] reg425 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg420 = (1'h0);
  reg [(4'h9):(1'h0)] reg419 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg417 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg416 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar412 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg411 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg410 = (1'h0);
  reg [(5'h12):(1'h0)] forvar407 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar406 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg403 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar402 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar395 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg394 = (1'h0);
  reg [(2'h2):(1'h0)] forvar393 = (1'h0);
  reg [(4'hc):(1'h0)] forvar391 = (1'h0);
  reg [(5'h13):(1'h0)] reg385 = (1'h0);
  reg [(5'h16):(1'h0)] reg389 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar388 = (1'h0);
  reg [(4'hc):(1'h0)] reg387 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg386 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar385 = (1'h0);
  reg [(2'h3):(1'h0)] reg384 = (1'h0);
  reg [(3'h5):(1'h0)] reg383 = (1'h0);
  reg [(5'h16):(1'h0)] reg382 = (1'h0);
  reg [(5'h18):(1'h0)] forvar381 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg380 = (1'h0);
  reg [(4'he):(1'h0)] forvar379 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg378 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg377 = (1'h0);
  reg [(4'hb):(1'h0)] reg375 = (1'h0);
  reg [(4'he):(1'h0)] reg374 = (1'h0);
  reg [(4'hb):(1'h0)] forvar369 = (1'h0);
  reg [(5'h16):(1'h0)] reg368 = (1'h0);
  reg [(5'h14):(1'h0)] reg367 = (1'h0);
  reg [(5'h17):(1'h0)] reg361 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg359 = (1'h0);
  reg [(4'h9):(1'h0)] reg358 = (1'h0);
  reg [(5'h16):(1'h0)] forvar357 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg356 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg355 = (1'h0);
  reg signed [(4'he):(1'h0)] reg354 = (1'h0);
  reg [(2'h2):(1'h0)] reg350 = (1'h0);
  reg [(4'hf):(1'h0)] reg348 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg347 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar344 = (1'h0);
  reg [(4'hf):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar341 = (1'h0);
  reg [(4'h9):(1'h0)] reg340 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg337 = (1'h0);
  reg [(4'hd):(1'h0)] reg335 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar333 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg332 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg331 = (1'h0);
  reg [(5'h12):(1'h0)] reg330 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg325 = (1'h0);
  reg [(2'h3):(1'h0)] reg328 = (1'h0);
  reg [(5'h14):(1'h0)] reg327 = (1'h0);
  reg [(5'h18):(1'h0)] forvar325 = (1'h0);
  reg [(3'h7):(1'h0)] reg321 = (1'h0);
  reg [(2'h3):(1'h0)] reg319 = (1'h0);
  reg [(4'he):(1'h0)] forvar318 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg317 = (1'h0);
  reg [(2'h2):(1'h0)] reg315 = (1'h0);
  reg [(5'h13):(1'h0)] reg314 = (1'h0);
  reg [(5'h17):(1'h0)] forvar313 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg311 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg309 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar307 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg305 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar301 = (1'h0);
  reg [(2'h3):(1'h0)] reg285 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg296 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg295 = (1'h0);
  reg [(5'h14):(1'h0)] reg294 = (1'h0);
  reg [(5'h12):(1'h0)] reg293 = (1'h0);
  reg [(3'h7):(1'h0)] reg291 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg290 = (1'h0);
  reg [(4'h9):(1'h0)] reg289 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg287 = (1'h0);
  reg [(2'h3):(1'h0)] reg286 = (1'h0);
  reg [(5'h10):(1'h0)] forvar285 = (1'h0);
  reg [(2'h2):(1'h0)] reg283 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg281 = (1'h0);
  reg [(5'h11):(1'h0)] reg279 = (1'h0);
  reg [(5'h17):(1'h0)] reg278 = (1'h0);
  reg [(4'hf):(1'h0)] forvar275 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg276 = (1'h0);
  reg [(4'hb):(1'h0)] reg274 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg272 = (1'h0);
  reg [(3'h6):(1'h0)] reg271 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg269 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg268 = (1'h0);
  reg [(5'h17):(1'h0)] reg265 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar264 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar261 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg259 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg258 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg255 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg252 = (1'h0);
  reg [(5'h11):(1'h0)] reg251 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg250 = (1'h0);
  reg [(4'hd):(1'h0)] reg246 = (1'h0);
  reg [(5'h14):(1'h0)] reg245 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg243 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg241 = (1'h0);
  reg [(3'h5):(1'h0)] forvar240 = (1'h0);
  reg [(4'h9):(1'h0)] reg239 = (1'h0);
  reg [(5'h10):(1'h0)] reg236 = (1'h0);
  reg [(5'h10):(1'h0)] reg235 = (1'h0);
  reg [(3'h7):(1'h0)] reg233 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg232 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg229 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg228 = (1'h0);
  reg [(5'h14):(1'h0)] reg222 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg220 = (1'h0);
  reg [(3'h6):(1'h0)] forvar219 = (1'h0);
  reg [(3'h5):(1'h0)] reg218 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg217 = (1'h0);
  reg [(4'hf):(1'h0)] forvar216 = (1'h0);
  reg [(5'h12):(1'h0)] reg215 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar213 = (1'h0);
  reg [(3'h4):(1'h0)] reg212 = (1'h0);
  reg [(3'h7):(1'h0)] forvar211 = (1'h0);
  reg [(5'h11):(1'h0)] reg209 = (1'h0);
  reg [(3'h5):(1'h0)] reg208 = (1'h0);
  reg [(4'h8):(1'h0)] reg207 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg206 = (1'h0);
  reg [(5'h18):(1'h0)] reg205 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg200 = (1'h0);
  assign y = {wire507,
                 wire424,
                 wire324,
                 wire249,
                 wire248,
                 wire247,
                 wire226,
                 wire225,
                 wire224,
                 reg490,
                 reg504,
                 reg502,
                 reg501,
                 reg496,
                 reg495,
                 reg493,
                 reg488,
                 reg485,
                 reg482,
                 reg481,
                 reg480,
                 reg476,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 reg469,
                 reg466,
                 reg460,
                 reg457,
                 reg456,
                 reg455,
                 reg453,
                 reg451,
                 reg450,
                 reg449,
                 reg447,
                 reg446,
                 reg441,
                 reg440,
                 reg438,
                 reg436,
                 reg435,
                 reg434,
                 reg432,
                 reg430,
                 reg428,
                 reg427,
                 reg426,
                 reg423,
                 reg422,
                 reg421,
                 reg418,
                 reg415,
                 reg413,
                 reg409,
                 reg408,
                 reg405,
                 reg404,
                 reg401,
                 reg400,
                 reg399,
                 reg398,
                 reg397,
                 reg396,
                 reg392,
                 reg390,
                 reg388,
                 reg376,
                 reg373,
                 reg372,
                 reg371,
                 reg370,
                 reg366,
                 reg365,
                 reg364,
                 reg363,
                 reg362,
                 reg360,
                 reg353,
                 reg352,
                 reg351,
                 reg349,
                 reg346,
                 reg345,
                 reg343,
                 reg342,
                 reg339,
                 reg338,
                 reg333,
                 reg336,
                 reg334,
                 reg329,
                 reg326,
                 reg313,
                 reg323,
                 reg322,
                 reg320,
                 reg316,
                 reg310,
                 reg307,
                 reg306,
                 reg304,
                 reg303,
                 reg302,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg292,
                 reg288,
                 reg284,
                 reg282,
                 reg280,
                 reg277,
                 reg275,
                 reg273,
                 reg270,
                 reg267,
                 reg266,
                 reg263,
                 reg262,
                 reg260,
                 reg257,
                 reg256,
                 reg254,
                 reg240,
                 reg244,
                 reg242,
                 reg238,
                 reg237,
                 reg234,
                 reg231,
                 reg230,
                 reg227,
                 reg223,
                 reg214,
                 reg210,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg497,
                 forvar496,
                 reg494,
                 forvar491,
                 reg506,
                 reg505,
                 forvar503,
                 reg500,
                 reg499,
                 reg498,
                 forvar497,
                 forvar494,
                 reg492,
                 reg491,
                 forvar490,
                 reg489,
                 reg487,
                 reg486,
                 reg484,
                 reg483,
                 reg479,
                 reg478,
                 forvar477,
                 reg475,
                 reg474,
                 reg468,
                 reg467,
                 reg465,
                 forvar452,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg459,
                 forvar458,
                 reg454,
                 reg452,
                 reg448,
                 forvar445,
                 reg444,
                 forvar443,
                 forvar442,
                 forvar434,
                 forvar425,
                 reg439,
                 reg437,
                 reg433,
                 reg431,
                 reg429,
                 reg425,
                 reg420,
                 reg419,
                 reg417,
                 reg416,
                 reg414,
                 forvar412,
                 reg411,
                 reg410,
                 forvar407,
                 forvar406,
                 reg403,
                 forvar402,
                 forvar395,
                 reg394,
                 forvar393,
                 forvar391,
                 reg385,
                 reg389,
                 forvar388,
                 reg387,
                 reg386,
                 forvar385,
                 reg384,
                 reg383,
                 reg382,
                 forvar381,
                 reg380,
                 forvar379,
                 reg378,
                 reg377,
                 reg375,
                 reg374,
                 forvar369,
                 reg368,
                 reg367,
                 reg361,
                 reg359,
                 reg358,
                 forvar357,
                 reg356,
                 reg355,
                 reg354,
                 reg350,
                 reg348,
                 reg347,
                 forvar344,
                 reg344,
                 forvar341,
                 reg340,
                 reg337,
                 reg335,
                 forvar333,
                 reg332,
                 reg331,
                 reg330,
                 reg325,
                 reg328,
                 reg327,
                 forvar325,
                 reg321,
                 reg319,
                 forvar318,
                 reg317,
                 reg315,
                 reg314,
                 forvar313,
                 reg312,
                 reg311,
                 reg309,
                 reg308,
                 forvar307,
                 reg305,
                 forvar301,
                 reg285,
                 reg296,
                 reg295,
                 reg294,
                 reg293,
                 reg291,
                 reg290,
                 reg289,
                 reg287,
                 reg286,
                 forvar285,
                 reg283,
                 reg281,
                 reg279,
                 reg278,
                 forvar275,
                 reg276,
                 reg274,
                 reg272,
                 reg271,
                 reg269,
                 reg268,
                 reg265,
                 forvar264,
                 forvar261,
                 reg259,
                 reg258,
                 reg255,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg246,
                 reg245,
                 reg243,
                 reg241,
                 forvar240,
                 reg239,
                 reg236,
                 reg235,
                 reg233,
                 reg232,
                 reg229,
                 reg228,
                 reg222,
                 reg221,
                 reg220,
                 forvar219,
                 reg218,
                 reg217,
                 forvar216,
                 reg215,
                 forvar213,
                 reg212,
                 forvar211,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg200,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((wire198 ?
          $signed(($unsigned($signed(wire199)) + ($unsigned(wire199) << {wire199,
              wire197}))) : wire196[(2'h3):(2'h2)]))
        begin
          reg200 = wire197;
          reg201 <= (((+{$signed(wire198)}) ?
                  (~((wire198 - wire199) ?
                      {wire198} : $signed(wire196))) : $signed(($unsigned(reg200) ?
                      $unsigned(wire198) : wire198))) ?
              ((((~|reg200) ? (reg200 ? wire199 : (7'h48)) : wire197) ?
                      wire197 : ((~&reg200) ?
                          {wire199, wire199} : $signed((8'ha7)))) ?
                  (-$unsigned(wire198)) : wire197) : $unsigned(wire197[(4'hd):(1'h0)]));
          reg202 <= ($unsigned((^~($unsigned(wire196) != (wire198 ?
              wire197 : wire196)))) << (-reg201));
          reg203 <= ((7'h4a) ?
              ($signed((!{wire196})) ?
                  reg200 : ({(wire197 | reg202)} ?
                      ({wire196} ^ (wire197 ?
                          wire196 : wire196)) : reg202)) : ({{wire198[(3'h7):(1'h1)]},
                  ($unsigned(wire199) && wire196[(4'he):(1'h0)])} - (~&$signed((~|(8'hbd))))));
          reg204 <= wire196;
        end
      else
        begin
          reg201 <= (+(wire197[(4'hd):(1'h0)] <= wire197[(4'hc):(4'h8)]));
          if ((reg202 > reg201[(2'h2):(1'h0)]))
            begin
              reg202 <= {(+$unsigned(wire196[(4'h8):(3'h5)])),
                  $unsigned((~&$unsigned(reg203[(3'h7):(3'h7)])))};
              reg203 <= (&({wire196[(4'h9):(4'h9)]} != $signed(reg204[(5'h15):(5'h12)])));
              reg205 = $unsigned($unsigned(({(~|wire199),
                  (wire196 ? wire199 : reg202)} >>> {$unsigned(reg201),
                  (reg201 ? reg202 : reg201)})));
            end
          else
            begin
              reg205 = $signed($unsigned(wire196));
              reg206 = {wire196};
              reg207 = $unsigned($unsigned(wire197[(4'ha):(1'h0)]));
              reg208 = $unsigned(wire198);
            end
          reg209 = (reg206 ? reg208 : reg205[(5'h13):(3'h4)]);
        end
      reg210 <= reg200;
      for (forvar211 = (1'h0); (forvar211 < (1'h0)); forvar211 = (forvar211 + (1'h1)))
        begin
          reg212 = (((|(&{reg200, (7'h45)})) ?
                  {$signed($unsigned(wire196)),
                      (~(7'h4a))} : $signed($signed(reg206))) ?
              reg210[(1'h0):(1'h0)] : (($unsigned($signed(wire199)) ^~ $signed(reg203)) || (($signed(reg202) ?
                      reg205 : $unsigned((8'hae))) ?
                  (8'ha9) : wire197[(3'h6):(1'h1)])));
          for (forvar213 = (1'h0); (forvar213 < (1'h0)); forvar213 = (forvar213 + (1'h1)))
            begin
              reg214 <= (~|($unsigned((^~$signed(wire196))) == ((~^$unsigned(reg202)) ?
                  reg206 : {(reg202 != wire199)})));
            end
          reg215 = reg214[(3'h4):(3'h4)];
        end
      for (forvar216 = (1'h0); (forvar216 < (2'h2)); forvar216 = (forvar216 + (1'h1)))
        begin
          reg217 = (!reg204);
          reg218 = ($signed((reg206 ?
              {(reg215 ?
                      forvar213 : (8'ha3))} : reg201)) & {(reg212[(1'h0):(1'h0)] ?
                  (^(reg207 ? reg212 : reg207)) : {(reg202 > wire197)})});
          for (forvar219 = (1'h0); (forvar219 < (3'h4)); forvar219 = (forvar219 + (1'h1)))
            begin
              reg220 = {((&(-(8'hb6))) ?
                      $signed(($signed(reg212) ?
                          $signed(forvar211) : {reg218,
                              reg203})) : (|((~^reg203) ?
                          $unsigned(reg208) : {reg200}))),
                  (8'hbe)};
              reg221 = {reg207[(1'h1):(1'h0)]};
              reg222 = $unsigned(($unsigned((reg218 - (reg202 ?
                      reg201 : wire196))) ?
                  reg204[(4'he):(4'hc)] : (reg207 || reg203)));
            end
        end
      reg223 <= $signed(reg209);
    end
  assign wire224 = reg202;
  assign wire225 = ({($unsigned($unsigned(reg223)) ?
                           $unsigned({reg223,
                               (8'h9d)}) : reg203[(4'hc):(3'h5)]),
                       reg223[(3'h6):(2'h3)]} > (((^~(~|reg223)) ?
                           wire197[(4'hb):(3'h6)] : $signed(reg204)) ?
                       reg214[(2'h3):(2'h2)] : $unsigned(($signed(reg204) && (reg202 ?
                           wire224 : wire224)))));
  assign wire226 = ($unsigned((((wire199 ? wire224 : reg214) ?
                           reg214 : wire224) ?
                       wire197 : $unsigned(reg203[(3'h4):(1'h1)]))) ^~ (($signed(reg204[(4'hd):(2'h2)]) ~^ {(reg223 + wire224)}) ?
                       $signed((&wire196[(3'h7):(1'h0)])) : $unsigned(reg214[(3'h4):(1'h1)])));
  always
    @(posedge clk) begin
      reg227 <= wire199[(1'h1):(1'h0)];
      reg228 = (~|reg227);
      if (((wire225[(4'hc):(2'h3)] >> reg201[(2'h2):(1'h1)]) ?
          (wire224 ?
              $signed($unsigned($unsigned((8'ha7)))) : (reg204[(4'hc):(3'h5)] >>> reg202[(3'h7):(3'h5)])) : {reg228[(3'h4):(3'h4)]}))
        begin
          if ($signed($signed($unsigned(reg223[(3'h4):(1'h1)]))))
            begin
              reg229 = reg202;
              reg230 <= reg210[(2'h3):(1'h1)];
            end
          else
            begin
              reg229 = $unsigned(reg228[(2'h2):(1'h1)]);
              reg230 <= wire224[(1'h1):(1'h1)];
              reg231 <= (wire224 ?
                  ({{(~&reg210)},
                          ((reg229 ? reg227 : reg203) * ((8'hae) - reg230))} ?
                      $unsigned(reg223[(3'h6):(1'h1)]) : ($unsigned($unsigned(reg227)) ?
                          (~reg229[(2'h2):(1'h0)]) : wire196[(4'hc):(2'h2)])) : ((((reg228 && reg228) && $signed(wire225)) && $unsigned(reg203[(1'h1):(1'h1)])) ?
                      (((!reg214) ?
                          (wire224 ?
                              wire196 : (7'h41)) : {wire197}) >>> $unsigned($signed(reg227))) : {$unsigned(reg230[(5'h16):(4'h9)])}));
            end
          if ($signed(reg214[(1'h1):(1'h0)]))
            begin
              reg232 = wire224[(4'h9):(2'h2)];
              reg233 = (-reg201[(3'h4):(3'h4)]);
              reg234 <= $signed(($signed($signed(wire199[(1'h1):(1'h0)])) ~^ reg210));
              reg235 = {$signed((&wire198[(3'h4):(2'h3)]))};
            end
          else
            begin
              reg234 <= $signed(reg230);
              reg235 = (~&$unsigned((({(8'hbf)} ?
                      wire198[(3'h5):(1'h1)] : $unsigned(wire198)) ?
                  $unsigned((wire226 | (8'ha6))) : ($unsigned(reg223) ^ (reg234 ?
                      reg231 : reg210)))));
              reg236 = reg233[(1'h1):(1'h1)];
              reg237 <= (~^$unsigned((wire197[(2'h3):(1'h0)] ?
                  (|(reg231 ^~ wire226)) : (reg204[(3'h5):(2'h2)] - (reg227 ~^ reg210)))));
              reg238 <= (~reg232[(2'h2):(1'h0)]);
            end
          reg239 = (8'ha6);
          for (forvar240 = (1'h0); (forvar240 < (3'h4)); forvar240 = (forvar240 + (1'h1)))
            begin
              reg241 = (($signed(reg223[(3'h6):(1'h0)]) ?
                      $signed(reg202) : {reg201[(1'h0):(1'h0)]}) ?
                  reg238[(1'h1):(1'h1)] : reg201);
              reg242 <= $signed((~&$signed(reg227)));
              reg243 = $unsigned(reg228[(2'h3):(1'h1)]);
              reg244 <= (($unsigned({(!forvar240)}) + $signed($signed((reg243 ?
                  reg243 : wire196)))) <= {$signed(($signed((8'hb5)) && ((8'had) ?
                      (8'hbe) : reg227)))});
              reg245 = ($signed(reg243) ?
                  wire198[(4'hc):(3'h6)] : ({((reg244 <= reg238) ?
                          (7'h48) : reg239[(3'h5):(1'h0)])} <<< reg223));
            end
          reg246 = $signed(reg242);
        end
      else
        begin
          reg229 = ((wire225[(1'h1):(1'h0)] ?
                  (8'hb5) : $unsigned({(wire196 ? (8'hbe) : reg233),
                      $signed(reg244)})) ?
              (reg233[(3'h4):(3'h4)] ?
                  reg237[(5'h14):(3'h4)] : $unsigned(reg238[(2'h3):(2'h2)])) : reg244);
          if (reg210)
            begin
              reg230 <= $signed($unsigned($unsigned(((reg231 ?
                  reg234 : (8'hb7)) << $signed(reg203)))));
              reg232 = $signed(forvar240[(1'h0):(1'h0)]);
              reg234 <= reg239;
            end
          else
            begin
              reg230 <= ($unsigned(reg202) >= reg241);
              reg232 = ((($signed((reg235 ^~ wire198)) && reg234) ?
                  wire199[(2'h3):(1'h0)] : {$unsigned((+reg243))}) + (~|wire224[(1'h0):(1'h0)]));
              reg234 <= reg234[(1'h1):(1'h1)];
            end
          reg237 <= reg233;
          reg239 = ((reg210 ?
              $signed(((|reg244) <<< {wire226})) : (~$signed(((7'h49) >>> reg204)))) <= ({{(8'hbd),
                      wire196[(3'h7):(3'h4)]}} ?
              ($signed(reg238) ?
                  $signed($signed(reg244)) : reg244[(3'h7):(1'h1)]) : $unsigned(reg228[(2'h3):(2'h2)])));
          reg240 <= ($signed(reg203) ?
              $unsigned(reg214[(3'h4):(1'h0)]) : $signed((8'had)));
        end
    end
  assign wire247 = {{($signed($signed(wire196)) ?
                               reg244[(1'h1):(1'h1)] : $signed((reg203 >>> reg201))),
                           ({$unsigned(wire224)} ?
                               $unsigned((reg202 ?
                                   reg240 : reg244)) : reg242[(4'ha):(4'h8)])}};
  assign wire248 = reg238;
  assign wire249 = $unsigned($signed(wire248[(4'ha):(2'h2)]));
  always
    @(posedge clk) begin
      reg250 = $signed({reg201[(2'h2):(1'h0)], reg214[(1'h0):(1'h0)]});
      reg251 = reg242[(4'hb):(2'h2)];
      if (((reg201[(3'h4):(2'h3)] * wire197) ?
          $signed((|(~|(reg250 ?
              reg210 : (7'h4a))))) : $unsigned({$unsigned($unsigned(reg230))})))
        begin
          reg252 = ((^(-(8'h9e))) ? (7'h41) : $unsigned(reg237));
          reg253 = $signed((~(((reg244 == reg214) >>> (wire225 - (8'h9d))) ?
              {((7'h41) ? wire224 : reg223),
                  $unsigned(reg238)} : (!(reg242 * reg230)))));
          reg254 <= (~&reg204[(5'h18):(4'hd)]);
          if ({($signed($signed(((8'hae) || (7'h49)))) == reg244[(4'ha):(1'h1)]),
              reg254})
            begin
              reg255 = (~|(8'hb9));
              reg256 <= reg201;
              reg257 <= (reg210 ?
                  $unsigned(wire247[(3'h5):(3'h4)]) : $signed($unsigned(reg251)));
            end
          else
            begin
              reg256 <= ({(reg210[(3'h7):(3'h7)] ?
                          $unsigned({reg227,
                              reg240}) : $signed($unsigned((7'h43))))} ?
                  $unsigned(reg231[(4'ha):(4'h8)]) : ($unsigned((wire199[(3'h6):(3'h6)] ?
                          $unsigned(wire198) : $signed(reg257))) ?
                      $unsigned(reg230[(4'hb):(3'h7)]) : $signed((8'ha7))));
              reg258 = reg234;
            end
          reg259 = (&($unsigned($signed({reg252})) ?
              wire199[(3'h7):(3'h4)] : (|$signed(wire247[(4'h8):(1'h0)]))));
        end
      else
        begin
          if ((8'hbd))
            begin
              reg252 = (reg258[(4'he):(2'h3)] ?
                  ((-wire247[(3'h7):(3'h6)]) >= (^~(8'hbb))) : reg244[(3'h6):(2'h3)]);
            end
          else
            begin
              reg252 = {$signed((-$signed(wire198))), wire247};
              reg253 = (7'h40);
            end
          if ((!reg242[(2'h2):(1'h0)]))
            begin
              reg254 <= reg227;
              reg255 = reg255[(5'h10):(3'h5)];
              reg256 <= wire248;
              reg257 <= (reg237 != (~|(({reg257, reg240} + (!reg254)) ?
                  reg257[(5'h13):(4'hc)] : $signed(reg230))));
              reg258 = $unsigned($signed((!(^$unsigned(reg234)))));
            end
          else
            begin
              reg255 = (((((reg255 ? reg237 : reg257) ?
                          $unsigned(wire198) : $signed(reg240)) ?
                      {reg252[(1'h0):(1'h0)]} : $unsigned($unsigned((8'hb2)))) + (8'haf)) ?
                  ($signed((|{reg251, wire197})) ?
                      {($unsigned(reg202) >>> (reg253 >>> wire249)),
                          (^~reg231)} : (((reg242 ?
                              (8'hb4) : reg253) >>> $signed(reg210)) ?
                          ($unsigned(reg240) ?
                              (wire225 <= (8'hb3)) : $unsigned(reg201)) : ((&(8'haa)) ?
                              wire198 : reg231))) : ($signed({reg255[(4'hd):(1'h1)],
                      reg238[(2'h3):(1'h1)]}) ^~ (^~(~^(reg227 ?
                      reg251 : reg210)))));
              reg258 = $signed((&reg259[(3'h4):(1'h1)]));
              reg260 <= (reg240 ?
                  $unsigned((((reg237 ? wire197 : wire199) ?
                          reg256 : $signed(reg251)) ?
                      $unsigned($unsigned(wire225)) : $signed((reg238 - reg257)))) : (wire198 || wire196));
            end
          for (forvar261 = (1'h0); (forvar261 < (1'h0)); forvar261 = (forvar261 + (1'h1)))
            begin
              reg262 <= reg238;
            end
          reg263 <= reg234[(1'h0):(1'h0)];
          for (forvar264 = (1'h0); (forvar264 < (1'h1)); forvar264 = (forvar264 + (1'h1)))
            begin
              reg265 = $signed(forvar264[(1'h1):(1'h0)]);
              reg266 <= (!$unsigned(reg204[(5'h18):(4'hb)]));
              reg267 <= ((~|({reg223[(4'h8):(1'h0)]} ?
                  ((wire196 ? reg253 : (8'ha7)) ?
                      (reg204 ?
                          reg214 : reg259) : (|reg244)) : (reg266[(5'h14):(4'hd)] * (reg237 ~^ reg257)))) - ({reg257[(4'h8):(3'h5)],
                      $signed((reg204 ? (8'hba) : forvar264))} ?
                  (!reg202[(3'h4):(1'h0)]) : wire197[(5'h10):(4'ha)]));
              reg268 = {(reg251[(4'hd):(3'h6)] * reg203)};
            end
        end
      reg269 = $unsigned(reg203[(4'hc):(3'h5)]);
      reg270 <= $unsigned(reg244[(4'h8):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg271 = $signed($signed($signed({{(8'ha9), (8'hb3)}, (|(8'hb5))})));
      if ((~$signed((^~$signed($unsigned(reg256))))))
        begin
          reg272 = {(($signed(wire224) ? reg234 : reg254) <<< (wire224 ?
                  (~(-(8'ha1))) : $signed((reg223 ? reg270 : reg227))))};
          if (({$signed(($unsigned(reg231) ? (!(8'haa)) : $unsigned(reg254)))} ?
              wire197[(4'h8):(3'h4)] : $unsigned(wire198)))
            begin
              reg273 <= $unsigned($signed(((^~reg271) ?
                  wire248[(1'h1):(1'h1)] : (8'ha0))));
              reg274 = ($unsigned(reg238) ? reg240[(4'h8):(1'h0)] : reg201);
            end
          else
            begin
              reg273 <= reg210[(2'h2):(1'h0)];
              reg275 <= (~reg242);
            end
          reg276 = (~$unsigned({(~^$unsigned((8'hae))),
              $unsigned((reg273 | reg274))}));
          reg277 <= reg271[(2'h3):(2'h3)];
        end
      else
        begin
          reg273 <= reg234;
          reg274 = (8'ha7);
          for (forvar275 = (1'h0); (forvar275 < (1'h1)); forvar275 = (forvar275 + (1'h1)))
            begin
              reg276 = reg277[(4'h8):(2'h2)];
              reg278 = (|(&(reg223[(2'h2):(1'h1)] == (8'ha0))));
            end
        end
      if (((wire198[(4'h9):(1'h1)] ?
          wire226 : reg204) == $signed({($signed(reg231) >= (reg262 << reg274)),
          $unsigned((7'h48))})))
        begin
          if (wire225[(1'h0):(1'h0)])
            begin
              reg279 = reg275;
              reg280 <= (({((^~reg223) ? (+reg214) : $signed(wire224)),
                          $unsigned(((8'ha6) ? reg256 : reg278))} ?
                      $unsigned(wire197) : ($unsigned((wire225 ?
                              reg210 : reg267)) ?
                          ((8'hb9) ?
                              reg278 : (reg203 ?
                                  reg262 : (7'h48))) : $signed((|reg277)))) ?
                  $unsigned($signed($unsigned((^reg271)))) : reg279);
              reg281 = (^~((-$unsigned((reg256 > reg244))) | (((~reg214) ?
                  {forvar275} : reg263[(2'h2):(2'h2)]) || wire226)));
              reg282 <= reg210;
              reg283 = (~^$unsigned({(reg234[(4'ha):(3'h5)] ?
                      (wire247 ? (7'h46) : reg231) : $unsigned(wire247))}));
            end
          else
            begin
              reg279 = ($signed((-reg223[(2'h2):(1'h1)])) ?
                  $unsigned((-reg267[(4'ha):(1'h0)])) : reg203[(3'h5):(1'h1)]);
              reg281 = (~|reg202);
              reg282 <= (~|$signed($signed(((reg279 - reg242) ?
                  reg280 : reg202))));
            end
          reg284 <= reg273;
          for (forvar285 = (1'h0); (forvar285 < (2'h2)); forvar285 = (forvar285 + (1'h1)))
            begin
              reg286 = ($unsigned({reg277[(2'h2):(1'h0)]}) ~^ $signed(($signed((reg284 != reg273)) ?
                  $signed($unsigned(reg278)) : reg276)));
              reg287 = reg237[(2'h3):(1'h0)];
              reg288 <= $signed($unsigned(reg231[(4'hb):(1'h1)]));
            end
          if ({{wire224}})
            begin
              reg289 = reg230[(3'h7):(2'h3)];
              reg290 = reg273;
              reg291 = ({$unsigned((^~$signed(reg201)))} ?
                  reg238 : $signed({$signed($unsigned(reg266))}));
            end
          else
            begin
              reg292 <= ($signed({$signed(((8'ha2) ?
                      reg237 : reg210))}) * wire224[(2'h2):(1'h0)]);
              reg293 = (~|(($signed((-reg267)) ?
                      wire198 : $signed((^~reg288))) ?
                  {$unsigned((wire226 ? (8'hab) : reg271))} : ((~reg263) ?
                      (8'h9d) : wire247[(4'hf):(1'h1)])));
              reg294 = (~^$signed((reg287[(4'ha):(4'h9)] < ((reg234 ?
                      reg267 : wire249) ?
                  reg281[(4'hf):(2'h2)] : $signed(reg257)))));
              reg295 = reg260;
              reg296 = ((8'ha0) ?
                  (wire196[(3'h6):(3'h5)] * wire196[(3'h6):(1'h0)]) : reg281[(2'h2):(1'h0)]);
            end
          reg297 <= (reg256[(4'hb):(1'h0)] && forvar285);
        end
      else
        begin
          if (wire198[(1'h1):(1'h0)])
            begin
              reg280 <= reg289[(3'h6):(2'h2)];
              reg281 = ((((reg280[(4'h8):(2'h3)] ~^ ((8'hb1) >= reg295)) ?
                      (((8'hab) ? reg280 : reg201) ?
                          ((7'h49) ? reg266 : reg271) : (reg280 ?
                              reg271 : reg223)) : reg291) != reg263) ?
                  wire196 : (&$signed($signed($unsigned(reg286)))));
              reg282 <= $signed((reg295[(3'h4):(2'h2)] || reg238));
              reg284 <= $unsigned(reg293);
              reg285 = (|((~reg242[(4'hb):(3'h5)]) ?
                  forvar285[(4'hf):(1'h0)] : ((8'hb8) ?
                      (reg286 ?
                          ((8'ha0) ?
                              reg230 : reg273) : reg223[(1'h0):(1'h0)]) : $signed($unsigned(reg295)))));
            end
          else
            begin
              reg279 = reg223[(3'h4):(3'h4)];
            end
          reg288 <= $unsigned(reg294);
          reg289 = (~^(reg201 < reg285));
          if ((reg202 - reg254[(3'h5):(1'h0)]))
            begin
              reg290 = reg254;
              reg292 <= $signed(forvar275);
              reg297 <= reg227[(1'h1):(1'h1)];
              reg298 <= (!reg203[(2'h2):(1'h1)]);
            end
          else
            begin
              reg292 <= ((reg231 ?
                      reg230[(3'h7):(3'h7)] : $signed($signed(reg227[(1'h0):(1'h0)]))) ?
                  (!$signed($unsigned((wire224 ?
                      reg257 : reg296)))) : $signed(($signed($signed(reg227)) & reg285[(1'h1):(1'h0)])));
              reg297 <= reg204;
              reg298 <= ((7'h44) - $unsigned((((~wire199) ? (8'hb0) : reg277) ?
                  ((forvar285 ? (7'h48) : reg201) ?
                      (wire198 ?
                          reg267 : (7'h4a)) : $signed(reg275)) : $unsigned(((8'ha8) ^~ reg279)))));
              reg299 <= $signed(wire199);
              reg300 <= reg267;
            end
          for (forvar301 = (1'h0); (forvar301 < (2'h3)); forvar301 = (forvar301 + (1'h1)))
            begin
              reg302 <= $unsigned(reg278[(5'h14):(4'h8)]);
              reg303 <= $signed($unsigned($signed($unsigned($unsigned(reg299)))));
              reg304 <= ($signed(reg266[(5'h15):(5'h14)]) ?
                  ((($unsigned(reg298) > (^~reg267)) | (reg283 + {forvar275})) - reg302[(1'h1):(1'h0)]) : {reg234,
                      $unsigned($signed((reg204 ? reg298 : (8'hb9))))});
              reg305 = reg284[(4'h9):(3'h4)];
              reg306 <= reg273[(3'h5):(2'h3)];
            end
        end
      if ($signed(reg288))
        begin
          reg307 <= ((^$unsigned((^(wire198 ? forvar275 : reg210)))) && reg237);
        end
      else
        begin
          for (forvar307 = (1'h0); (forvar307 < (2'h3)); forvar307 = (forvar307 + (1'h1)))
            begin
              reg308 = reg214;
              reg309 = $signed((((&wire248[(2'h3):(1'h1)]) <= $unsigned((reg266 & reg256))) ?
                  $unsigned((((8'hb2) ? (8'h9f) : reg290) ?
                      (reg237 * (8'ha1)) : $unsigned(reg298))) : (|$unsigned((~^reg283)))));
              reg310 <= $signed($signed($unsigned($unsigned((reg227 ?
                  reg238 : reg308)))));
              reg311 = (-$unsigned(reg293[(4'hc):(4'h9)]));
            end
        end
      if (((7'h44) || wire226[(5'h14):(5'h10)]))
        begin
          reg312 = (+((7'h47) ?
              ($signed($unsigned(reg204)) ^~ (forvar275 ?
                  {reg242} : reg293[(4'hb):(3'h6)])) : {(+(|reg287)),
                  (-(wire248 ^~ reg273))}));
          for (forvar313 = (1'h0); (forvar313 < (1'h0)); forvar313 = (forvar313 + (1'h1)))
            begin
              reg314 = $unsigned($signed((reg296[(2'h2):(1'h0)] && $unsigned((reg262 <<< forvar307)))));
              reg315 = ((reg280[(3'h6):(1'h0)] ?
                      $signed({(^~wire226),
                          $unsigned(reg289)}) : $signed(reg308)) ?
                  (reg210 <<< reg285[(1'h1):(1'h0)]) : ((reg280[(2'h2):(1'h1)] ?
                      (reg286[(1'h1):(1'h0)] ?
                          reg297[(5'h13):(5'h13)] : $unsigned(forvar301)) : reg273) * $signed(((reg289 <= reg284) ?
                      (reg310 ? reg270 : reg298) : $signed(wire197)))));
              reg316 <= $unsigned(($signed($unsigned((|reg262))) ?
                  (reg298[(2'h3):(1'h0)] ?
                      (~^reg297[(5'h12):(4'hc)]) : ((wire225 ^ (7'h41)) * reg273[(4'h8):(1'h1)])) : wire224));
            end
          reg317 = $unsigned((^((-$unsigned(wire247)) < (|$unsigned(reg242)))));
          for (forvar318 = (1'h0); (forvar318 < (2'h2)); forvar318 = (forvar318 + (1'h1)))
            begin
              reg319 = (~&(!$unsigned(($signed((8'ha6)) || reg310))));
              reg320 <= $signed((~(reg305[(1'h0):(1'h0)] ^~ reg317[(1'h1):(1'h0)])));
              reg321 = {(+reg204),
                  $signed(($signed(reg237[(1'h1):(1'h0)]) != $signed((forvar313 | reg214))))};
              reg322 <= (|$signed({((reg300 ? forvar275 : reg311) ?
                      (reg291 ? reg320 : reg234) : $unsigned((7'h44)))}));
              reg323 <= (reg286 < (reg267[(2'h2):(1'h0)] ?
                  $signed(((reg312 ?
                      reg271 : reg280) << reg262[(4'hf):(4'hd)])) : {(~|reg296)}));
            end
        end
      else
        begin
          reg313 <= $signed($signed(($unsigned((reg202 ? wire249 : (8'hae))) ?
              ((reg278 ^~ reg321) ?
                  (reg234 ?
                      forvar301 : (7'h4a)) : reg322[(1'h1):(1'h0)]) : $signed((reg297 | (8'ha8))))));
          reg314 = {reg283[(2'h2):(2'h2)]};
        end
    end
  assign wire324 = {(((^~$signed(reg254)) ?
                           {$unsigned((8'hb8)), reg230} : ((reg288 ?
                               reg316 : reg234) == (^reg275))) ^ $unsigned($unsigned({reg201,
                           reg302})))};
  always
    @(posedge clk) begin
      if ($signed($unsigned(reg313)))
        begin
          for (forvar325 = (1'h0); (forvar325 < (2'h3)); forvar325 = (forvar325 + (1'h1)))
            begin
              reg326 <= (reg240[(4'h9):(4'h9)] ?
                  (~wire249) : (~$unsigned(reg273[(1'h1):(1'h0)])));
              reg327 = {((&$signed(reg298[(1'h1):(1'h1)])) >= (((reg260 ?
                              reg280 : reg275) ?
                          wire225 : reg302[(3'h7):(1'h0)]) ?
                      (|$signed(reg227)) : ((reg298 <<< reg299) ?
                          reg326 : wire249)))};
            end
          reg328 = reg323;
        end
      else
        begin
          reg325 = (~^wire248[(5'h10):(4'hd)]);
          if (reg323[(1'h1):(1'h0)])
            begin
              reg327 = (wire224[(3'h4):(1'h0)] ? $unsigned(reg300) : reg260);
            end
          else
            begin
              reg327 = $unsigned((-reg262));
              reg329 <= $unsigned(wire197);
              reg330 = (($signed((8'h9d)) ~^ ((((8'hb1) | (8'haa)) != $unsigned((7'h47))) ?
                  (reg304[(1'h1):(1'h0)] ?
                      reg325 : {reg273,
                          reg240}) : reg254)) > reg256[(5'h16):(4'h9)]);
              reg331 = reg242[(2'h3):(2'h2)];
              reg332 = (^($unsigned(((reg230 ~^ reg288) > $signed(wire198))) ?
                  reg282 : (~^reg227[(1'h1):(1'h0)])));
            end
        end
      if ((reg214 ? wire247[(4'hb):(1'h0)] : reg299[(4'hb):(4'hb)]))
        begin
          for (forvar333 = (1'h0); (forvar333 < (3'h4)); forvar333 = (forvar333 + (1'h1)))
            begin
              reg334 <= wire198[(1'h1):(1'h1)];
            end
          if (reg203)
            begin
              reg335 = (($signed(($unsigned(reg332) ?
                          $signed(reg316) : reg242[(4'h9):(1'h1)])) ?
                      ($unsigned($signed(reg238)) ?
                          reg280 : (!reg326)) : reg330) ?
                  wire248 : ($unsigned((((8'hb9) <= reg322) ?
                      (reg331 ?
                          reg334 : reg288) : $signed(reg304))) - (&{(reg242 ?
                          reg210 : wire324)})));
              reg336 <= ($unsigned($unsigned(({reg262,
                      reg325} >= (wire324 || reg335)))) ?
                  $signed(reg288[(4'he):(3'h7)]) : ((({reg330} ?
                      wire198 : (8'hba)) && $signed({reg238,
                      reg240})) << (reg256 ?
                      reg277[(3'h6):(3'h4)] : ($signed(reg304) == ((8'ha8) == (8'hbf))))));
            end
          else
            begin
              reg336 <= $signed($signed((((~|(8'had)) ?
                      reg275[(4'ha):(3'h4)] : $unsigned((8'ha7))) ?
                  reg304[(2'h2):(1'h1)] : (^reg277))));
            end
        end
      else
        begin
          if (reg227)
            begin
              reg333 <= wire247;
              reg334 <= $unsigned($unsigned($unsigned((^reg273[(3'h5):(2'h2)]))));
              reg336 <= wire324;
            end
          else
            begin
              reg335 = (((reg284[(5'h11):(1'h1)] >>> $unsigned(forvar325)) >> wire226[(5'h13):(3'h7)]) * $unsigned(reg262[(3'h5):(2'h3)]));
              reg336 <= reg307;
              reg337 = reg313;
            end
          reg338 <= {$unsigned((!((wire224 >> reg297) > (reg227 != reg302)))),
              $signed((-reg302[(3'h5):(1'h0)]))};
          if ((+($unsigned($unsigned($signed(reg329))) ?
              {$unsigned({reg273, wire248}),
                  $signed(wire248[(4'he):(4'hd)])} : (&(reg284[(4'hf):(1'h0)] ?
                  $signed(reg302) : $signed(reg303))))))
            begin
              reg339 <= $unsigned((reg320 - reg292));
              reg340 = {((8'ha5) && $signed((^$signed(reg275))))};
            end
          else
            begin
              reg339 <= reg223[(3'h6):(1'h1)];
              reg340 = reg339;
            end
          for (forvar341 = (1'h0); (forvar341 < (3'h4)); forvar341 = (forvar341 + (1'h1)))
            begin
              reg342 <= (~reg322[(3'h4):(2'h2)]);
              reg343 <= (~&($unsigned($unsigned(wire196[(4'he):(4'hb)])) == {reg332[(2'h3):(1'h1)],
                  wire225}));
            end
        end
      if (($signed(((!(reg297 ? reg335 : (7'h47))) ?
          wire199[(2'h2):(1'h0)] : reg282)) ^~ ((~$unsigned((reg334 ?
              reg298 : wire247))) ?
          (reg323 ?
              ($signed(reg306) ~^ (reg299 ? reg202 : reg288)) : {{reg322,
                      reg242},
                  $unsigned(reg322)}) : $signed(($signed(reg263) ?
              reg327[(3'h7):(3'h4)] : (reg300 + reg273))))))
        begin
          reg344 = (!{$unsigned(reg329[(4'he):(4'ha)])});
        end
      else
        begin
          for (forvar344 = (1'h0); (forvar344 < (1'h0)); forvar344 = (forvar344 + (1'h1)))
            begin
              reg345 <= reg302;
              reg346 <= reg310[(3'h4):(2'h3)];
              reg347 = reg334[(3'h7):(3'h6)];
            end
          reg348 = $signed((reg203 ?
              $unsigned($unsigned(reg331)) : ($unsigned(wire196[(5'h10):(4'hf)]) == (reg323[(4'h9):(1'h1)] ?
                  (-reg288) : (&reg242)))));
          if ((-reg325))
            begin
              reg349 <= (^~{(~reg347), reg270});
              reg350 = (8'hb0);
            end
          else
            begin
              reg349 <= (-(~^(reg292 ?
                  reg230[(4'ha):(2'h3)] : {$unsigned(reg275),
                      forvar333[(2'h2):(2'h2)]})));
              reg351 <= $unsigned(reg280[(2'h3):(2'h2)]);
              reg352 <= reg275;
            end
          reg353 <= (($unsigned(reg352[(2'h2):(1'h0)]) ?
              $unsigned(reg350) : $signed({reg302[(1'h0):(1'h0)]})) ^ (reg352 ?
              (-($signed((8'hb1)) ?
                  reg329[(3'h5):(1'h0)] : (~|reg307))) : reg327[(4'hb):(3'h5)]));
          reg354 = $unsigned({(reg323 ? reg227 : $unsigned($signed(reg254))),
              ($unsigned((reg336 ? wire248 : wire248)) ~^ forvar341)});
        end
      reg355 = (reg322 ?
          $unsigned($signed(((reg340 ? reg306 : wire197) ?
              (8'ha1) : $unsigned(reg322)))) : $signed({({reg203} ~^ ((8'hae) ?
                  (8'hac) : wire249))}));
    end
  always
    @(posedge clk) begin
      reg356 = ($unsigned(reg322[(3'h4):(1'h1)]) ?
          reg260 : $signed(((reg307[(2'h2):(2'h2)] ?
              reg320 : reg333[(1'h0):(1'h0)]) >> wire248)));
      for (forvar357 = (1'h0); (forvar357 < (3'h4)); forvar357 = (forvar357 + (1'h1)))
        begin
          if ($signed(((((~|(8'hb2)) || reg304) ?
                  (~|$signed(reg242)) : ((reg356 != reg263) ?
                      (reg270 <= reg275) : $signed((7'h43)))) ?
              $signed(((reg313 >>> reg277) ?
                  (~^reg234) : (~|reg300))) : ((!{(8'hba)}) ?
                  $unsigned((reg230 ? reg316 : reg257)) : reg201))))
            begin
              reg358 = (($signed(((reg203 ?
                      (8'had) : reg202) | $signed(reg214))) & $unsigned(((-reg223) ?
                      (+reg304) : $signed(reg353)))) ?
                  $unsigned(({$unsigned((8'h9c))} ?
                      reg260 : reg260[(1'h1):(1'h0)])) : reg231);
              reg359 = $signed($unsigned(reg298[(2'h3):(1'h0)]));
              reg360 <= reg227[(1'h0):(1'h0)];
              reg361 = (reg302 >> $signed($signed(($unsigned(reg351) ?
                  (|(8'hb7)) : (reg343 ? reg313 : wire198)))));
            end
          else
            begin
              reg360 <= reg284;
              reg361 = $signed(reg257[(5'h14):(4'he)]);
              reg362 <= reg356;
            end
          reg363 <= reg362;
          if (reg282[(5'h11):(4'hc)])
            begin
              reg364 <= reg266[(5'h10):(5'h10)];
              reg365 <= (+wire196[(3'h5):(1'h0)]);
              reg366 <= reg338;
            end
          else
            begin
              reg364 <= reg323;
              reg367 = (reg273[(2'h3):(2'h3)] ?
                  wire198[(4'hb):(2'h2)] : (!reg363));
              reg368 = ($unsigned({reg204}) && $signed(reg292[(1'h1):(1'h1)]));
            end
          for (forvar369 = (1'h0); (forvar369 < (1'h0)); forvar369 = (forvar369 + (1'h1)))
            begin
              reg370 <= reg302[(3'h7):(3'h7)];
            end
          if (($signed((reg234 ?
              (7'h46) : {wire198,
                  wire226[(4'hc):(4'hc)]})) <= wire248[(4'h8):(3'h4)]))
            begin
              reg371 <= $unsigned($unsigned(reg234));
              reg372 <= $unsigned($unsigned(wire197));
              reg373 <= wire324;
            end
          else
            begin
              reg371 <= $unsigned(((!$unsigned((reg349 ? reg371 : reg202))) ?
                  reg343[(1'h1):(1'h1)] : $signed((+reg203))));
              reg372 <= (reg227[(1'h1):(1'h0)] ?
                  $unsigned((((reg372 ? wire224 : reg204) >= (~|wire198)) ?
                      reg359[(1'h0):(1'h0)] : $unsigned(reg345[(2'h2):(2'h2)]))) : $signed(((!(reg275 > reg326)) >> $signed(wire324[(3'h7):(3'h7)]))));
              reg374 = (!((7'h43) ? $signed((!$signed(reg254))) : (|reg333)));
              reg375 = (reg334[(1'h0):(1'h0)] == (8'ha6));
              reg376 <= {(reg375[(1'h1):(1'h1)] <= (~|(((8'hac) ~^ wire197) ?
                      $unsigned(reg362) : $signed(reg343)))),
                  reg288};
            end
        end
    end
  always
    @(posedge clk) begin
      reg377 = ({$signed((reg310[(1'h1):(1'h1)] == reg353[(4'hc):(4'hc)])),
          (^(^~(reg333 ?
              reg376 : wire198)))} != (reg201[(2'h2):(1'h0)] ^ reg277));
    end
  always
    @(posedge clk) begin
      reg378 = (wire247 | (($unsigned($unsigned(reg240)) >>> reg284[(4'h8):(2'h2)]) <= $unsigned($signed($unsigned(reg336)))));
      for (forvar379 = (1'h0); (forvar379 < (1'h0)); forvar379 = (forvar379 + (1'h1)))
        begin
          reg380 = $signed(wire198);
          for (forvar381 = (1'h0); (forvar381 < (1'h0)); forvar381 = (forvar381 + (1'h1)))
            begin
              reg382 = ({(7'h4a), reg282[(5'h10):(1'h0)]} ?
                  reg339 : {$signed((~&$unsigned(reg302)))});
              reg383 = reg300;
            end
          reg384 = reg376[(4'h8):(3'h4)];
        end
      if ({reg304[(1'h0):(1'h0)]})
        begin
          for (forvar385 = (1'h0); (forvar385 < (3'h4)); forvar385 = (forvar385 + (1'h1)))
            begin
              reg386 = reg210;
              reg387 = (+reg310);
            end
          for (forvar388 = (1'h0); (forvar388 < (2'h3)); forvar388 = (forvar388 + (1'h1)))
            begin
              reg389 = (((8'h9f) ?
                      reg336[(3'h6):(1'h0)] : (^~(reg240 ? reg334 : reg288))) ?
                  reg370[(3'h4):(3'h4)] : (reg297 ?
                      forvar388[(1'h0):(1'h0)] : $unsigned(reg238[(2'h3):(1'h1)])));
            end
        end
      else
        begin
          if ((!reg345))
            begin
              reg385 = $unsigned((reg386 ~^ (+$unsigned($unsigned(reg223)))));
              reg388 <= $signed((reg256[(4'ha):(2'h2)] ?
                  (($signed((8'ha5)) < (reg389 ?
                      reg339 : reg364)) >>> (~(^reg242))) : reg227[(1'h0):(1'h0)]));
              reg390 <= (~(+forvar385[(3'h6):(1'h0)]));
            end
          else
            begin
              reg388 <= ((~(reg343[(4'hb):(4'hb)] >= (reg214 & {reg388}))) ?
                  (|(reg389 && $unsigned((7'h4a)))) : reg371[(4'hf):(4'hf)]);
              reg389 = $unsigned(((+((^~wire248) <<< $signed((8'ha7)))) ^ (^~(reg263[(3'h4):(2'h3)] ?
                  (+(7'h42)) : (7'h46)))));
            end
          for (forvar391 = (1'h0); (forvar391 < (3'h4)); forvar391 = (forvar391 + (1'h1)))
            begin
              reg392 <= (~|$signed({{$unsigned(reg372)}}));
            end
          for (forvar393 = (1'h0); (forvar393 < (2'h3)); forvar393 = (forvar393 + (1'h1)))
            begin
              reg394 = ($signed((8'hb6)) ?
                  ($unsigned(reg342) && ({$unsigned(reg223),
                          (reg388 < (8'haa))} ?
                      {forvar388[(4'hc):(1'h1)],
                          (reg204 ? (8'h9e) : reg366)} : ((reg360 ?
                          reg257 : reg284) | (wire248 - reg346)))) : $unsigned(($unsigned($signed(wire197)) ~^ forvar379[(4'h9):(3'h6)])));
            end
          for (forvar395 = (1'h0); (forvar395 < (2'h2)); forvar395 = (forvar395 + (1'h1)))
            begin
              reg396 <= {$unsigned(reg320), $signed(reg302)};
              reg397 <= $unsigned(reg302[(4'h9):(2'h2)]);
              reg398 <= (&reg353[(4'hd):(3'h5)]);
              reg399 <= reg244;
              reg400 <= {reg306};
            end
          reg401 <= reg380[(1'h0):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar402 = (1'h0); (forvar402 < (1'h1)); forvar402 = (forvar402 + (1'h1)))
        begin
          reg403 = $signed($signed({(^~(reg343 ? reg234 : reg397))}));
          reg404 <= (~|reg338);
          reg405 <= (reg353 | reg303);
        end
    end
  always
    @(posedge clk) begin
      for (forvar406 = (1'h0); (forvar406 < (3'h4)); forvar406 = (forvar406 + (1'h1)))
        begin
          for (forvar407 = (1'h0); (forvar407 < (3'h4)); forvar407 = (forvar407 + (1'h1)))
            begin
              reg408 <= (((^~reg282) != $unsigned(reg362[(1'h1):(1'h0)])) > forvar406);
              reg409 <= $unsigned(reg365[(1'h1):(1'h0)]);
              reg410 = (|(reg302 ?
                  $unsigned(reg234) : (~{reg304[(3'h5):(2'h3)]})));
            end
          reg411 = $unsigned(reg360);
          for (forvar412 = (1'h0); (forvar412 < (2'h2)); forvar412 = (forvar412 + (1'h1)))
            begin
              reg413 <= {(^~$unsigned((-$unsigned(reg270))))};
              reg414 = forvar412[(3'h6):(2'h2)];
            end
          if ((~|(reg336[(4'h8):(2'h3)] - wire249)))
            begin
              reg415 <= (wire249[(4'hf):(4'h9)] ?
                  (~^(wire247[(2'h3):(1'h1)] ?
                      (reg371 >>> (reg292 ?
                          reg256 : (8'had))) : wire249)) : ((|($unsigned(reg313) ?
                          (reg345 >>> reg345) : reg313)) ?
                      $signed($unsigned((reg256 ?
                          wire199 : reg376))) : reg297[(2'h3):(2'h3)]));
              reg416 = ({reg300[(1'h1):(1'h1)],
                      $signed(((wire197 ?
                          reg214 : reg297) == reg415[(4'ha):(3'h7)]))} ?
                  $unsigned($unsigned($unsigned((wire247 >> reg300)))) : $signed({(~&$unsigned(reg339)),
                      $signed(reg227[(1'h0):(1'h0)])}));
              reg417 = wire249[(4'ha):(3'h7)];
              reg418 <= reg352[(1'h0):(1'h0)];
            end
          else
            begin
              reg415 <= (reg204 != $unsigned($unsigned(((reg298 && wire324) >>> reg316))));
              reg416 = {($signed(reg342[(1'h1):(1'h1)]) > $signed((^~$signed(reg204)))),
                  (|$unsigned($signed(wire249)))};
              reg418 <= (7'h45);
              reg419 = $signed(reg376);
              reg420 = reg313[(3'h4):(1'h0)];
            end
        end
      reg421 <= $unsigned(reg323);
      reg422 <= $unsigned(reg322[(3'h6):(1'h1)]);
      reg423 <= $signed($signed((reg336 + ((reg292 ?
          reg338 : reg238) >>> reg409))));
    end
  assign wire424 = (7'h48);
  always
    @(posedge clk) begin
      if (((($unsigned(reg422) ?
              {reg257[(5'h10):(1'h1)]} : reg322[(1'h0):(1'h0)]) ?
          ({(reg401 || reg262), (reg423 * reg409)} <= ({reg349} ?
              wire324 : reg310)) : $signed({(reg342 ?
                  (8'hae) : wire197)})) ^ reg270))
        begin
          if ((~&reg231))
            begin
              reg425 = reg275;
              reg426 <= reg338;
              reg427 <= $unsigned($unsigned(((reg280[(3'h6):(1'h0)] ?
                      (7'h43) : (!reg266)) ?
                  $unsigned($unsigned(reg202)) : {((8'haa) >> reg320)})));
              reg428 <= (($signed($signed((8'ha2))) < $signed((reg230 & (wire248 * reg415)))) ?
                  $unsigned((({reg396} > $unsigned(reg298)) ?
                      $unsigned({reg363}) : reg282)) : $signed($signed($signed($signed(reg333)))));
            end
          else
            begin
              reg426 <= ((reg266 ^ ($signed($unsigned(reg349)) ?
                      ((reg401 >= reg310) < $signed(reg364)) : reg256)) ?
                  (~{$unsigned((!wire198)),
                      ((reg339 ? reg376 : wire199) ?
                          reg349 : (reg204 ? (8'hab) : reg313))}) : (8'hac));
              reg427 <= (+(~&(~|((~&reg277) ~^ (reg338 >> reg238)))));
              reg429 = (8'hba);
            end
          reg430 <= ($signed((reg373 << $signed((|reg345)))) ?
              {(|(8'hac))} : $signed(($signed($signed(reg231)) ?
                  {reg334[(4'h8):(1'h1)],
                      reg399[(1'h1):(1'h1)]} : {$unsigned(wire247)})));
          if (wire199)
            begin
              reg431 = (+{reg334[(4'hf):(1'h0)]});
              reg432 <= reg399;
              reg433 = $unsigned($unsigned($signed((~^reg306))));
            end
          else
            begin
              reg432 <= reg428;
            end
          reg434 <= $unsigned((~(((&reg234) | reg316[(5'h10):(3'h4)]) + $unsigned($unsigned(reg404)))));
          if ($unsigned(($signed((!((8'ha1) ? reg298 : wire226))) ~^ reg345)))
            begin
              reg435 <= ($unsigned($signed(({reg338,
                  reg280} < $signed(reg202)))) <<< ($unsigned({(reg399 >= reg346),
                  {reg307, reg262}}) >>> $signed($signed($unsigned(reg353)))));
              reg436 <= reg408[(2'h3):(1'h0)];
              reg437 = {reg282[(4'h8):(2'h2)],
                  $signed(($signed((reg390 == reg230)) != {(8'ha1),
                      $unsigned(reg362)}))};
              reg438 <= reg426[(2'h3):(1'h1)];
              reg439 = $unsigned((~^$signed({reg302, (7'h41)})));
            end
          else
            begin
              reg437 = ((reg388 ?
                  (-$signed(reg257[(4'hf):(4'hf)])) : reg244) >>> (reg244[(3'h4):(2'h2)] && $unsigned((&(~|(8'hbc))))));
              reg438 <= $unsigned(($unsigned((~$signed(reg203))) ?
                  {$unsigned($signed(reg277))} : wire196));
              reg440 <= reg421[(4'hd):(2'h3)];
              reg441 <= $unsigned({$signed(((~^wire324) ?
                      ((8'hb1) ? reg365 : reg298) : $unsigned(reg260)))});
            end
        end
      else
        begin
          for (forvar425 = (1'h0); (forvar425 < (2'h3)); forvar425 = (forvar425 + (1'h1)))
            begin
              reg426 <= reg438;
              reg427 <= reg303;
            end
          if ($signed(reg363[(1'h1):(1'h0)]))
            begin
              reg428 <= (&(reg372[(5'h13):(5'h12)] ?
                  $unsigned({(8'h9e),
                      (~|forvar425)}) : ((~&(&(7'h45))) >> $signed((reg415 ?
                      wire249 : reg320)))));
              reg430 <= (($signed(({reg339} | (^reg339))) ?
                  (((reg303 << reg345) ? $signed(reg431) : $signed(reg266)) ?
                      reg292[(2'h2):(1'h1)] : (reg421 >= (reg343 ?
                          (8'had) : reg254))) : reg428) >= (~|{(reg398 ?
                      reg423[(3'h6):(3'h5)] : reg231)}));
            end
          else
            begin
              reg429 = $unsigned($signed(({$unsigned((8'hae))} ?
                  reg254[(3'h6):(1'h0)] : $signed((|reg210)))));
              reg431 = (+(reg270 ?
                  $signed($signed((-reg282))) : {reg342[(4'h8):(1'h0)]}));
              reg432 <= ((reg415[(4'ha):(2'h3)] - (~$signed($unsigned(reg349)))) ?
                  reg263 : reg418[(1'h1):(1'h0)]);
              reg433 = (($unsigned(reg373) + wire424) ?
                  (|reg441[(3'h4):(1'h1)]) : $unsigned(($unsigned(reg343) >> reg282)));
            end
          for (forvar434 = (1'h0); (forvar434 < (3'h4)); forvar434 = (forvar434 + (1'h1)))
            begin
              reg435 <= $signed($signed((8'hb6)));
            end
        end
      for (forvar442 = (1'h0); (forvar442 < (2'h2)); forvar442 = (forvar442 + (1'h1)))
        begin
          for (forvar443 = (1'h0); (forvar443 < (2'h2)); forvar443 = (forvar443 + (1'h1)))
            begin
              reg444 = {reg349[(4'hf):(4'h9)]};
            end
          for (forvar445 = (1'h0); (forvar445 < (1'h0)); forvar445 = (forvar445 + (1'h1)))
            begin
              reg446 <= reg390[(3'h5):(2'h2)];
            end
        end
    end
  always
    @(posedge clk) begin
      if ((7'h4a))
        begin
          if (($signed((wire247[(4'he):(4'hc)] & (^~$signed(reg320)))) == reg326))
            begin
              reg447 <= $signed($signed($signed($signed($signed(reg322)))));
            end
          else
            begin
              reg448 = reg298;
              reg449 <= (($unsigned(reg345[(4'ha):(1'h0)]) ?
                      (+$unsigned((!reg427))) : ((~reg362[(3'h5):(1'h0)]) ?
                          $signed((8'hb6)) : $unsigned($unsigned(reg300)))) ?
                  (($signed(((7'h45) && reg204)) ?
                          reg202 : (reg401 >= reg320)) ?
                      (&{reg415[(3'h7):(3'h4)]}) : (reg427 & (&$signed((8'hba))))) : reg370);
              reg450 <= reg421;
            end
          if (($signed(reg441) <= {$unsigned($unsigned(((8'ha4) + reg307))),
              reg298[(2'h2):(1'h1)]}))
            begin
              reg451 <= $unsigned($unsigned($unsigned($signed(reg299[(4'he):(1'h1)]))));
              reg452 = {($signed(reg398[(4'hd):(4'h8)]) ?
                      reg440 : (~|(&(-reg263)))),
                  {reg430}};
              reg453 <= ({reg320} ?
                  wire196[(3'h5):(3'h5)] : ((reg427 * reg280[(1'h1):(1'h0)]) ?
                      reg435 : reg333));
              reg454 = $unsigned($signed((8'hbf)));
            end
          else
            begin
              reg451 <= wire424;
              reg453 <= reg371;
              reg455 <= $unsigned(({$signed(wire249[(4'hf):(4'hd)]),
                  (&{reg353, reg399})} != (((!(8'hba)) || (-reg438)) ?
                  (reg299 ?
                      reg275[(4'hf):(4'h8)] : {wire197,
                          reg275}) : $signed(((8'hb4) | reg436)))));
              reg456 <= $signed(({$signed((wire424 <<< reg333))} ?
                  ($unsigned(reg257) ^~ reg422) : reg342));
              reg457 <= reg204[(5'h11):(4'he)];
            end
          for (forvar458 = (1'h0); (forvar458 < (2'h2)); forvar458 = (forvar458 + (1'h1)))
            begin
              reg459 = reg423;
              reg460 <= reg435[(2'h3):(1'h0)];
              reg461 = (($signed($signed((~|reg231))) + reg438) ?
                  reg326[(4'hb):(4'hb)] : ({($signed(reg292) >> (reg396 + reg413)),
                          $signed((reg342 >> reg303))} ?
                      reg284[(4'hf):(3'h5)] : $unsigned($signed(((7'h4a) - reg267)))));
              reg462 = reg404[(4'he):(3'h5)];
              reg463 = $unsigned({($unsigned(reg329) >> ((&reg415) ?
                      (reg280 >> reg388) : $signed(reg397)))});
            end
          reg464 = reg266[(2'h3):(2'h2)];
        end
      else
        begin
          if ((wire249 >>> {reg260[(4'h9):(2'h3)]}))
            begin
              reg448 = ((~|reg310) ?
                  $unsigned(wire196) : ((^~reg372) || (~^$unsigned({reg300}))));
              reg449 <= {{(((reg397 ?
                          reg310 : (8'ha6)) << $unsigned((8'hb4))) >> {(!reg464),
                          {reg300}}),
                      (((reg223 < wire247) ?
                              $signed(reg292) : $unsigned(reg267)) ?
                          (&$signed(reg326)) : ({reg448} + (reg306 ~^ reg230)))}};
            end
          else
            begin
              reg447 <= $unsigned(reg460[(4'ha):(2'h2)]);
              reg449 <= {(-wire198), $signed(reg304[(3'h5):(1'h1)])};
              reg450 <= (forvar458[(1'h1):(1'h0)] && $signed(reg323[(1'h0):(1'h0)]));
              reg451 <= ($signed((reg238[(4'hd):(4'hb)] * (-reg427))) ?
                  $signed(reg270[(1'h0):(1'h0)]) : reg238[(4'h8):(1'h1)]);
            end
          for (forvar452 = (1'h0); (forvar452 < (2'h2)); forvar452 = (forvar452 + (1'h1)))
            begin
              reg454 = (&((((|wire224) * (reg204 ? reg460 : reg307)) ?
                  $signed((~^reg242)) : ($signed(reg422) * $unsigned((8'hbc)))) <= ($unsigned((!reg304)) ?
                  (8'hb8) : ((reg227 & reg349) > (reg398 ? reg370 : reg447)))));
              reg455 <= $unsigned($unsigned(reg438[(2'h3):(2'h2)]));
              reg456 <= reg455[(1'h0):(1'h0)];
            end
          reg457 <= ($signed($signed(reg202)) ? (~&reg339) : reg461);
        end
      if (reg388[(1'h0):(1'h0)])
        begin
          if ({$signed(reg201)})
            begin
              reg465 = (~((((8'h9f) ? reg463 : reg418) ?
                  ({reg288, reg242} | (~^reg266)) : ((~&reg434) ?
                      (&reg298) : reg270[(3'h5):(1'h1)])) <<< {(wire224 ?
                      $signed(reg257) : (!reg266))}));
              reg466 <= ((~&$signed({$signed(reg303)})) ?
                  reg237 : $unsigned((+$unsigned($unsigned((8'hbf))))));
              reg467 = ((7'h49) >= ((&reg297) >> (((~reg210) * {reg362}) | $signed((reg454 ?
                  reg401 : reg430)))));
              reg468 = (-reg303[(2'h3):(1'h1)]);
            end
          else
            begin
              reg465 = reg399;
              reg466 <= reg238[(4'h9):(4'h9)];
              reg469 <= reg418;
              reg470 <= reg401[(1'h0):(1'h0)];
              reg471 <= $signed($unsigned($signed(((forvar458 >> reg300) >= (reg307 ?
                  reg460 : reg303)))));
            end
          reg472 <= {wire324[(1'h0):(1'h0)], reg405};
          if ((+reg405[(3'h7):(3'h7)]))
            begin
              reg473 <= $signed({(^wire199), $unsigned((~|$signed(reg448)))});
              reg474 = reg273;
              reg475 = (reg323 ?
                  (^~reg352[(2'h3):(1'h1)]) : reg418[(3'h6):(3'h4)]);
            end
          else
            begin
              reg473 <= ($unsigned(reg396[(1'h1):(1'h1)]) ?
                  reg426[(1'h1):(1'h1)] : $unsigned({$unsigned(((8'ha0) ?
                          reg201 : reg254))}));
            end
        end
      else
        begin
          reg466 <= reg373[(3'h5):(2'h2)];
          if (reg430)
            begin
              reg469 <= $unsigned((((~^(reg298 ? (8'hb9) : reg360)) ?
                      reg201[(1'h1):(1'h0)] : {(~&reg372)}) ?
                  $unsigned((((8'haa) ? reg270 : reg351) ?
                      reg470[(5'h12):(4'hb)] : (~&(8'hb0)))) : $signed((((8'hb8) ?
                          reg463 : reg227) ?
                      (reg467 & reg230) : (8'h9e)))));
              reg474 = $unsigned(reg284[(4'h9):(3'h6)]);
              reg476 <= ($unsigned((reg300[(2'h2):(2'h2)] ?
                      $signed($unsigned(reg280)) : $unsigned(((8'hbc) ?
                          reg447 : reg372)))) ?
                  reg438[(1'h1):(1'h1)] : ((((!reg364) ?
                              (~|wire424) : ((8'hb2) ? wire197 : reg462)) ?
                          $unsigned((~|reg270)) : reg202) ?
                      $signed(reg267) : $unsigned((8'hbe))));
            end
          else
            begin
              reg467 = $signed((reg365 && (~&$unsigned($signed(wire224)))));
              reg468 = reg376;
              reg469 <= reg299;
            end
          for (forvar477 = (1'h0); (forvar477 < (2'h2)); forvar477 = (forvar477 + (1'h1)))
            begin
              reg478 = $unsigned((|(8'hb2)));
              reg479 = (!reg447[(1'h1):(1'h1)]);
              reg480 <= (|($unsigned(reg401[(3'h5):(3'h4)]) <= $unsigned(reg415)));
            end
          reg481 <= ($unsigned(((reg260[(2'h2):(2'h2)] ?
                  (reg292 ? reg370 : reg334) : reg474[(1'h0):(1'h0)]) ?
              (~$unsigned(reg455)) : $unsigned(reg456))) < $signed(({(wire324 ?
                      reg460 : reg392),
                  $unsigned(wire225)} ?
              $unsigned(wire247) : (~|$signed(reg244)))));
        end
      if (reg464)
        begin
          if ($signed((+(reg202 ?
              reg426 : ({reg333, reg260} ?
                  $signed(reg336) : $unsigned(reg409))))))
            begin
              reg482 <= reg303[(1'h1):(1'h0)];
              reg483 = reg475[(5'h12):(4'hd)];
              reg484 = ($signed((~|reg449[(4'ha):(1'h0)])) ?
                  {reg464[(1'h1):(1'h1)],
                      $unsigned(reg388[(1'h1):(1'h1)])} : $unsigned($unsigned(($unsigned(reg231) ?
                      $unsigned(reg362) : (reg376 == reg364)))));
              reg485 <= {reg474,
                  ((~&$signed((reg483 ? reg329 : reg277))) ?
                      reg329[(3'h4):(1'h1)] : (($signed(reg326) ?
                              (^~reg310) : {reg202}) ?
                          reg277[(4'h8):(3'h6)] : reg284[(5'h13):(4'hf)]))};
            end
          else
            begin
              reg483 = (((!wire249[(5'h14):(3'h6)]) ?
                      $signed(((wire249 <= reg453) > ((7'h42) + reg399))) : ($unsigned((reg234 ?
                          (7'h49) : wire198)) >>> ((reg363 ?
                          (8'hbb) : reg303) <<< (reg450 == reg320)))) ?
                  {(reg460[(1'h0):(1'h0)] ?
                          ({reg366} ?
                              (reg397 ? reg470 : (8'ha9)) : (reg413 ?
                                  reg430 : reg244)) : ((-reg352) <<< (|reg237)))} : $unsigned($unsigned($signed((reg334 & (8'ha8))))));
              reg485 <= $signed(reg260[(5'h13):(4'he)]);
              reg486 = reg468[(4'hc):(3'h6)];
              reg487 = $signed(($unsigned($signed((reg481 <<< reg408))) ?
                  $unsigned(wire249) : (8'haa)));
              reg488 <= (({(reg270[(2'h3):(2'h2)] ?
                          reg462 : $signed(reg364))} && ($unsigned(reg284) ?
                      ($signed(reg326) || $unsigned(reg400)) : (((7'h47) ?
                          reg203 : wire324) >> $unsigned((8'had))))) ?
                  (7'h41) : ($signed($signed((^reg478))) ?
                      (^~{(reg303 ~^ reg484)}) : $signed(((!reg266) ?
                          (reg446 < reg487) : {reg409, reg418}))));
            end
        end
      else
        begin
          if (((~&reg409) ?
              {reg455,
                  ($unsigned((reg428 ?
                      reg487 : reg322)) - $unsigned(((8'ha7) <<< reg275)))} : (^(reg426[(3'h5):(1'h1)] ^ $unsigned((reg464 ?
                  reg413 : reg455))))))
            begin
              reg483 = reg413;
            end
          else
            begin
              reg483 = reg468;
            end
          reg485 <= (~|reg334[(4'h9):(2'h2)]);
          reg488 <= ($unsigned((&(~|$signed(reg237)))) ?
              {((~^((7'h47) ? reg399 : reg427)) << ((~(7'h48)) ?
                      {reg430, (7'h44)} : $signed(reg257))),
                  reg413[(3'h5):(1'h0)]} : $unsigned($signed(($signed(reg435) ?
                  {reg392, reg353} : (^reg401)))));
        end
      reg489 = $unsigned($signed(($unsigned(reg284) != ((reg334 ^ reg452) >> (reg230 ?
          (8'hb0) : (8'hab))))));
      if (reg352)
        begin
          for (forvar490 = (1'h0); (forvar490 < (2'h3)); forvar490 = (forvar490 + (1'h1)))
            begin
              reg491 = (^$unsigned($unsigned((^~(~&reg436)))));
              reg492 = ((~|((reg363[(2'h2):(2'h2)] ?
                      reg203 : reg478[(4'h9):(3'h4)]) ?
                  $signed({(8'hbb),
                      reg372}) : (reg478 & (^~reg302)))) == reg488);
              reg493 <= reg320;
            end
          for (forvar494 = (1'h0); (forvar494 < (1'h1)); forvar494 = (forvar494 + (1'h1)))
            begin
              reg495 <= ($unsigned(($unsigned((^~reg326)) ^ (8'haf))) >>> (~^($signed(reg288) ?
                  {$unsigned(wire199), {reg434, reg334}} : reg452)));
              reg496 <= (~{(8'hb0), {reg365}});
            end
          for (forvar497 = (1'h0); (forvar497 < (2'h2)); forvar497 = (forvar497 + (1'h1)))
            begin
              reg498 = ((reg280 || ($unsigned(reg299[(1'h1):(1'h0)]) ?
                      ($signed(reg238) ?
                          $unsigned(reg334) : reg316[(3'h5):(1'h1)]) : (reg404 != (^reg485)))) ?
                  reg440 : $unsigned((&(~(^reg365)))));
              reg499 = ($unsigned((-$signed((reg364 ? reg310 : (8'had))))) ?
                  ((+({(7'h49)} ? (reg496 ? wire224 : reg352) : (&reg320))) ?
                      $signed(reg441[(1'h1):(1'h0)]) : (!reg313)) : $unsigned(($signed((wire248 ?
                          reg459 : reg365)) ?
                      (+(reg400 == wire424)) : reg426[(1'h1):(1'h0)])));
              reg500 = reg453[(5'h17):(3'h5)];
              reg501 <= reg496;
            end
          reg502 <= {(reg404[(4'hd):(3'h4)] && $signed($signed(reg446))),
              wire197[(5'h10):(4'hc)]};
          for (forvar503 = (1'h0); (forvar503 < (1'h1)); forvar503 = (forvar503 + (1'h1)))
            begin
              reg504 <= reg351[(2'h2):(1'h1)];
              reg505 = reg447;
              reg506 = $unsigned($unsigned((reg300[(1'h1):(1'h0)] ?
                  {reg434} : {(~|reg491), ((8'had) ? reg282 : reg408)})));
            end
        end
      else
        begin
          reg490 <= reg266;
          for (forvar491 = (1'h0); (forvar491 < (3'h4)); forvar491 = (forvar491 + (1'h1)))
            begin
              reg492 = reg490;
              reg494 = (+(({(reg475 ? reg371 : wire196), $unsigned(forvar477)} ?
                  (|(^reg326)) : $unsigned(wire199)) != (~&reg342)));
              reg495 <= ((reg397 ?
                      $signed($unsigned($signed(reg476))) : (($signed(reg388) ?
                          reg502[(2'h2):(2'h2)] : $unsigned(reg316)) <<< $unsigned($signed(reg405)))) ?
                  $unsigned({$unsigned((reg210 >> reg254)),
                      {reg434[(2'h3):(1'h0)]}}) : $signed(reg489[(4'h9):(1'h1)]));
            end
          for (forvar496 = (1'h0); (forvar496 < (3'h4)); forvar496 = (forvar496 + (1'h1)))
            begin
              reg497 = {(reg237[(5'h14):(5'h10)] ?
                      (((reg485 >> reg266) <= (reg336 ?
                          reg481 : reg464)) < $unsigned(reg469)) : {$unsigned($signed((7'h49)))}),
                  (-(reg496 ?
                      ((reg473 ? reg326 : reg284) ?
                          (~&reg415) : ((7'h43) ?
                              reg292 : reg451)) : ((reg470 && (8'hba)) ^ reg362[(4'ha):(1'h0)])))};
              reg498 = ($unsigned($signed(reg473)) & $unsigned({$signed((8'hb7)),
                  $unsigned($signed((8'h9f)))}));
              reg499 = reg487[(3'h4):(2'h3)];
            end
          reg501 <= $signed({reg421[(5'h13):(5'h10)]});
        end
    end
  assign wire507 = (8'haa);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1432
#(parameter param1592 = {(({((8'hb2) ? (8'ha4) : (7'h42)), ((8'h9e) ? (8'hba) : (8'hb5))} ? (((8'ha5) ? (8'hba) : (7'h48)) ? (^(8'hb4)) : ((8'haa) ? (8'had) : (8'hb3))) : ((^(8'hb0)) ? ((8'hb3) >> (8'hbd)) : ((8'ha8) + (8'hb3)))) ? (!(((8'hbb) == (8'h9c)) - ((7'h43) ~^ (8'hab)))) : ((((8'ha6) ? (8'hbb) : (8'hb7)) ? (!(8'ha5)) : ((8'h9d) ? (8'haa) : (8'hb3))) == (((8'ha2) || (8'hbf)) ? ((8'hb4) ^~ (7'h4a)) : (-(8'haa)))))})
(y, clk, wire1436, wire1435, wire1434, wire1433);
  output wire [(32'h86c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire1436;
  input wire [(4'he):(1'h0)] wire1435;
  input wire [(4'hc):(1'h0)] wire1434;
  input wire signed [(5'h10):(1'h0)] wire1433;
  wire signed [(4'ha):(1'h0)] wire1564;
  wire [(4'ha):(1'h0)] wire1563;
  wire [(5'h13):(1'h0)] wire1523;
  wire signed [(5'h13):(1'h0)] wire1522;
  wire [(4'hd):(1'h0)] wire1521;
  wire signed [(2'h3):(1'h0)] wire1480;
  wire signed [(4'hf):(1'h0)] wire1479;
  wire [(5'h15):(1'h0)] wire1465;
  wire signed [(5'h16):(1'h0)] wire1464;
  wire [(3'h6):(1'h0)] wire1453;
  reg signed [(5'h11):(1'h0)] reg1588 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1580 = (1'h0);
  reg [(3'h5):(1'h0)] reg1579 = (1'h0);
  reg [(4'he):(1'h0)] reg1578 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1577 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1574 = (1'h0);
  reg [(5'h14):(1'h0)] reg1567 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1561 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1557 = (1'h0);
  reg [(5'h18):(1'h0)] reg1553 = (1'h0);
  reg [(3'h4):(1'h0)] reg1558 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1556 = (1'h0);
  reg [(4'hd):(1'h0)] reg1554 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1551 = (1'h0);
  reg [(4'hf):(1'h0)] reg1549 = (1'h0);
  reg [(4'h8):(1'h0)] reg1548 = (1'h0);
  reg [(4'hd):(1'h0)] reg1547 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1545 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1542 = (1'h0);
  reg [(4'he):(1'h0)] reg1541 = (1'h0);
  reg [(5'h10):(1'h0)] reg1538 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1535 = (1'h0);
  reg [(5'h14):(1'h0)] reg1533 = (1'h0);
  reg [(5'h12):(1'h0)] reg1532 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1530 = (1'h0);
  reg [(4'he):(1'h0)] reg1528 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1527 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1526 = (1'h0);
  reg [(4'hf):(1'h0)] reg1524 = (1'h0);
  reg [(4'hd):(1'h0)] reg1519 = (1'h0);
  reg [(4'he):(1'h0)] reg1514 = (1'h0);
  reg [(2'h3):(1'h0)] reg1513 = (1'h0);
  reg [(5'h13):(1'h0)] reg1510 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1508 = (1'h0);
  reg [(4'h9):(1'h0)] reg1507 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1506 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1502 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1501 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1498 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1496 = (1'h0);
  reg [(5'h12):(1'h0)] reg1495 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1494 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1493 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1490 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1486 = (1'h0);
  reg [(5'h10):(1'h0)] reg1485 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1476 = (1'h0);
  reg [(4'ha):(1'h0)] reg1475 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1460 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1458 = (1'h0);
  reg [(3'h4):(1'h0)] reg1457 = (1'h0);
  reg [(4'ha):(1'h0)] reg1456 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1450 = (1'h0);
  reg [(3'h5):(1'h0)] reg1448 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1445 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1443 = (1'h0);
  reg [(4'hb):(1'h0)] reg1442 = (1'h0);
  reg [(5'h11):(1'h0)] reg1441 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1440 = (1'h0);
  reg [(5'h11):(1'h0)] reg1439 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1438 = (1'h0);
  reg [(5'h13):(1'h0)] reg1437 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1591 = (1'h0);
  reg [(4'hb):(1'h0)] reg1590 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1589 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1587 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1586 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1585 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1584 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1583 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1582 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1581 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1576 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1575 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1573 = (1'h0);
  reg [(5'h11):(1'h0)] reg1572 = (1'h0);
  reg [(3'h5):(1'h0)] reg1571 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1570 = (1'h0);
  reg [(4'he):(1'h0)] reg1569 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1568 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1566 = (1'h0);
  reg [(4'he):(1'h0)] reg1565 = (1'h0);
  reg [(5'h17):(1'h0)] reg1562 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1556 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1551 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1546 = (1'h0);
  reg [(4'hd):(1'h0)] reg1560 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1559 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1557 = (1'h0);
  reg [(5'h13):(1'h0)] reg1555 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar1553 = (1'h0);
  reg [(5'h14):(1'h0)] reg1552 = (1'h0);
  reg [(3'h7):(1'h0)] reg1550 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1546 = (1'h0);
  reg [(5'h10):(1'h0)] reg1544 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1543 = (1'h0);
  reg [(4'h8):(1'h0)] reg1540 = (1'h0);
  reg [(4'hf):(1'h0)] reg1539 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1537 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1536 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1534 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1530 = (1'h0);
  reg [(3'h4):(1'h0)] reg1529 = (1'h0);
  reg [(4'hd):(1'h0)] reg1531 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1529 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1525 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1520 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1518 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1517 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1516 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1515 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1512 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1511 = (1'h0);
  reg [(4'ha):(1'h0)] reg1509 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1505 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1504 = (1'h0);
  reg [(3'h4):(1'h0)] reg1503 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1500 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1499 = (1'h0);
  reg [(5'h14):(1'h0)] reg1497 = (1'h0);
  reg [(5'h18):(1'h0)] reg1492 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1491 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1489 = (1'h0);
  reg [(5'h18):(1'h0)] reg1488 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1484 = (1'h0);
  reg [(5'h16):(1'h0)] reg1487 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1484 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1483 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1482 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1481 = (1'h0);
  reg [(5'h17):(1'h0)] reg1478 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1477 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1474 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1473 = (1'h0);
  reg [(3'h6):(1'h0)] reg1472 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1471 = (1'h0);
  reg [(2'h2):(1'h0)] reg1470 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1469 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1468 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1467 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1466 = (1'h0);
  reg [(3'h5):(1'h0)] reg1463 = (1'h0);
  reg [(5'h18):(1'h0)] reg1462 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1461 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1459 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1455 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1454 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1452 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1451 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1449 = (1'h0);
  reg [(4'hc):(1'h0)] reg1447 = (1'h0);
  reg [(4'hc):(1'h0)] reg1446 = (1'h0);
  reg [(4'hb):(1'h0)] reg1444 = (1'h0);
  assign y = {wire1564,
                 wire1563,
                 wire1523,
                 wire1522,
                 wire1521,
                 wire1480,
                 wire1479,
                 wire1465,
                 wire1464,
                 wire1453,
                 reg1588,
                 reg1580,
                 reg1579,
                 reg1578,
                 reg1577,
                 reg1574,
                 reg1567,
                 reg1561,
                 reg1557,
                 reg1553,
                 reg1558,
                 reg1556,
                 reg1554,
                 reg1551,
                 reg1549,
                 reg1548,
                 reg1547,
                 reg1545,
                 reg1542,
                 reg1541,
                 reg1538,
                 reg1535,
                 reg1533,
                 reg1532,
                 reg1530,
                 reg1528,
                 reg1527,
                 reg1526,
                 reg1524,
                 reg1519,
                 reg1514,
                 reg1513,
                 reg1510,
                 reg1508,
                 reg1507,
                 reg1506,
                 reg1502,
                 reg1501,
                 reg1498,
                 reg1496,
                 reg1495,
                 reg1494,
                 reg1493,
                 reg1490,
                 reg1486,
                 reg1485,
                 reg1476,
                 reg1475,
                 reg1460,
                 reg1458,
                 reg1457,
                 reg1456,
                 reg1450,
                 reg1448,
                 reg1445,
                 reg1443,
                 reg1442,
                 reg1441,
                 reg1440,
                 reg1439,
                 reg1438,
                 reg1437,
                 reg1591,
                 reg1590,
                 reg1589,
                 forvar1587,
                 reg1586,
                 reg1585,
                 reg1584,
                 reg1583,
                 reg1582,
                 forvar1581,
                 reg1576,
                 reg1575,
                 reg1573,
                 reg1572,
                 reg1571,
                 reg1570,
                 reg1569,
                 reg1568,
                 reg1566,
                 reg1565,
                 reg1562,
                 forvar1556,
                 forvar1551,
                 forvar1546,
                 reg1560,
                 reg1559,
                 forvar1557,
                 reg1555,
                 forvar1553,
                 reg1552,
                 reg1550,
                 reg1546,
                 reg1544,
                 reg1543,
                 reg1540,
                 reg1539,
                 forvar1537,
                 reg1536,
                 reg1534,
                 forvar1530,
                 reg1529,
                 reg1531,
                 forvar1529,
                 forvar1525,
                 reg1520,
                 forvar1518,
                 reg1517,
                 reg1516,
                 forvar1515,
                 reg1512,
                 reg1511,
                 reg1509,
                 reg1505,
                 forvar1504,
                 reg1503,
                 reg1500,
                 reg1499,
                 reg1497,
                 reg1492,
                 reg1491,
                 reg1489,
                 reg1488,
                 reg1484,
                 reg1487,
                 forvar1484,
                 reg1483,
                 reg1482,
                 reg1481,
                 reg1478,
                 reg1477,
                 reg1474,
                 reg1473,
                 reg1472,
                 reg1471,
                 reg1470,
                 reg1469,
                 reg1468,
                 reg1467,
                 forvar1466,
                 reg1463,
                 reg1462,
                 reg1461,
                 reg1459,
                 reg1455,
                 forvar1454,
                 reg1452,
                 reg1451,
                 reg1449,
                 reg1447,
                 reg1446,
                 reg1444,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1437 <= (($unsigned((wire1434 == $signed(wire1433))) | wire1435[(3'h4):(2'h3)]) ?
          ($unsigned(wire1434[(2'h3):(2'h2)]) << ((~^{wire1433,
              wire1434}) >= (^(~^wire1433)))) : wire1436[(4'he):(4'ha)]);
      if ((-$signed(reg1437[(4'he):(2'h2)])))
        begin
          reg1438 <= ($unsigned($unsigned((!$unsigned(reg1437)))) > {(^((wire1434 - (8'hbf)) && $signed(wire1433))),
              (reg1437[(5'h12):(4'h8)] * wire1434)});
        end
      else
        begin
          if ((7'h48))
            begin
              reg1438 <= ($unsigned((~^(wire1434[(4'hc):(4'h8)] ?
                      reg1437[(3'h6):(3'h6)] : $unsigned(wire1436)))) ?
                  ((wire1436[(3'h7):(2'h3)] * (~^(wire1435 ?
                      wire1436 : wire1435))) ~^ $unsigned(wire1433)) : $unsigned((wire1434 != $unsigned((wire1434 != (8'hbd))))));
              reg1439 <= ({(((wire1434 ? reg1437 : reg1438) ?
                      $unsigned(wire1435) : ((8'hb7) >>> reg1438)) != ($signed(wire1433) == (wire1436 ?
                      reg1437 : wire1433)))} & wire1434[(4'h8):(2'h2)]);
              reg1440 <= (-(~wire1435));
              reg1441 <= (((|($signed(reg1437) ?
                      wire1433[(4'hd):(3'h5)] : (~|reg1439))) ?
                  $signed((reg1437 ?
                      $unsigned(wire1436) : $unsigned((8'h9d)))) : reg1439) >= $unsigned((~^(-reg1440))));
            end
          else
            begin
              reg1438 <= $signed($unsigned((~&((-reg1438) & wire1436[(3'h7):(3'h4)]))));
            end
        end
      if (reg1441[(1'h1):(1'h0)])
        begin
          reg1442 <= (|wire1433[(3'h4):(2'h2)]);
          reg1443 <= $unsigned((!($signed((reg1442 || wire1434)) + $signed($signed(wire1436)))));
          reg1444 = {$signed({wire1434, ((8'hbf) & {wire1435})}),
              (wire1433[(4'h9):(3'h7)] >= ((-(wire1435 ~^ (8'hbf))) ^ $signed($signed(reg1443))))};
          reg1445 <= ({{reg1439,
                  ($signed((8'hb5)) ~^ $unsigned(wire1434))}} ~^ reg1443[(4'h9):(1'h0)]);
        end
      else
        begin
          reg1444 = $signed({(({reg1444} ? (8'hb9) : {reg1437}) || (reg1438 ?
                  $signed(reg1443) : reg1442))});
          if ((reg1440[(2'h3):(1'h0)] ?
              reg1445 : ($unsigned((8'ha6)) ?
                  $signed((^((7'h48) ?
                      reg1443 : wire1434))) : {{(reg1445 << wire1433),
                          (reg1445 ? reg1438 : reg1444)}})))
            begin
              reg1446 = (~($unsigned(($signed(wire1433) ?
                      reg1444[(2'h2):(1'h0)] : $signed(reg1440))) ?
                  {$unsigned((~|reg1444)),
                      reg1438[(2'h2):(2'h2)]} : (({reg1445} ?
                          wire1433[(4'he):(4'h8)] : (reg1438 ?
                              reg1439 : (8'hb0))) ?
                      {$signed((7'h48))} : reg1442[(1'h1):(1'h1)])));
              reg1447 = (+($signed(reg1439) >= (~|(-$signed(reg1437)))));
              reg1448 <= reg1444[(2'h2):(1'h0)];
              reg1449 = reg1448;
              reg1450 <= reg1443;
            end
          else
            begin
              reg1445 <= $unsigned(((~|{{reg1437}}) ?
                  $unsigned((-(reg1448 ? (8'hbe) : (7'h45)))) : wire1434));
              reg1448 <= reg1447[(1'h0):(1'h0)];
              reg1449 = $unsigned(wire1433);
            end
          reg1451 = $signed(wire1435);
        end
      reg1452 = {reg1448[(1'h1):(1'h1)]};
    end
  assign wire1453 = $signed((^reg1437));
  always
    @(posedge clk) begin
      for (forvar1454 = (1'h0); (forvar1454 < (2'h3)); forvar1454 = (forvar1454 + (1'h1)))
        begin
          reg1455 = $unsigned(wire1435[(4'he):(2'h3)]);
          reg1456 <= ((8'hb8) ? reg1455 : reg1437);
          reg1457 <= wire1453;
          reg1458 <= $unsigned((^($signed(wire1434[(1'h0):(1'h0)]) - $unsigned($unsigned(reg1455)))));
          reg1459 = reg1437;
        end
      reg1460 <= forvar1454[(3'h7):(2'h2)];
      reg1461 = reg1448;
      reg1462 = reg1461[(3'h7):(1'h0)];
      reg1463 = ($unsigned({$unsigned({reg1459, reg1448}),
              {$signed(wire1434)}}) ?
          ($unsigned((^~$signed(wire1436))) >= {wire1435[(3'h5):(2'h2)],
              $unsigned((wire1434 ?
                  reg1462 : reg1450))}) : $signed($signed(reg1443[(3'h7):(1'h0)])));
    end
  assign wire1464 = $unsigned((reg1450 * reg1440[(4'he):(4'he)]));
  assign wire1465 = (~&wire1433[(4'hc):(3'h4)]);
  always
    @(posedge clk) begin
      for (forvar1466 = (1'h0); (forvar1466 < (2'h2)); forvar1466 = (forvar1466 + (1'h1)))
        begin
          if (($unsigned($unsigned((~reg1448))) >>> ($unsigned($unsigned(reg1450[(3'h4):(3'h4)])) ?
              {$unsigned(reg1438[(2'h2):(2'h2)])} : $unsigned(((8'hbc) ?
                  (reg1437 ? (8'hb5) : reg1460) : (~&(8'hbe)))))))
            begin
              reg1467 = $signed((reg1443[(4'ha):(1'h0)] ?
                  wire1434 : reg1441[(4'he):(2'h2)]));
              reg1468 = ($unsigned(reg1450[(4'h8):(3'h4)]) && $signed(reg1438[(1'h0):(1'h0)]));
              reg1469 = (($unsigned(reg1460[(2'h3):(2'h2)]) ?
                  $signed((&(reg1458 | reg1439))) : $signed($unsigned({reg1445,
                      (8'hbc)}))) && (8'ha4));
            end
          else
            begin
              reg1467 = wire1433[(4'h9):(3'h7)];
            end
          if ($unsigned($unsigned((($unsigned(reg1457) ^ $signed((8'hb9))) ?
              (^reg1450[(4'hc):(3'h5)]) : reg1437[(4'h8):(3'h4)]))))
            begin
              reg1470 = $signed($signed($signed(wire1436[(3'h7):(1'h1)])));
              reg1471 = $signed(((($unsigned(reg1468) ?
                      wire1434[(3'h7):(1'h1)] : reg1458[(2'h2):(1'h1)]) >>> $signed(wire1464)) ?
                  $unsigned($unsigned((~reg1440))) : $unsigned({wire1433[(4'h9):(3'h6)],
                      {reg1440, (7'h4a)}})));
              reg1472 = {reg1469};
              reg1473 = (((forvar1466[(3'h7):(3'h4)] <<< $unsigned((~|(8'ha0)))) ^~ ((~&$signed(wire1433)) && {(reg1471 ?
                      wire1464 : wire1436)})) + reg1438[(3'h5):(3'h5)]);
              reg1474 = ($unsigned(wire1464) ~^ ($unsigned(reg1441[(4'h8):(2'h2)]) ^ $signed($unsigned(reg1458))));
            end
          else
            begin
              reg1470 = (~&reg1445);
              reg1475 <= (-$signed((($unsigned(reg1441) ?
                      $unsigned((7'h42)) : $unsigned((8'hbd))) ?
                  {{wire1433, reg1439}} : $unsigned({reg1448}))));
              reg1476 <= (((~&reg1467) ?
                  {($unsigned(reg1439) || (reg1468 && (8'hbe))),
                      ((reg1458 > (7'h4a)) ?
                          {reg1456} : (reg1468 ?
                              reg1469 : (8'hb6)))} : $unsigned(((wire1464 < reg1468) <<< wire1465[(4'he):(3'h7)]))) <= (($signed($signed(wire1453)) ?
                  $unsigned((~&reg1445)) : (reg1474 ?
                      (7'h4a) : $unsigned(wire1436))) <<< ({(&reg1458)} | reg1467[(3'h7):(1'h0)])));
              reg1477 = reg1439;
              reg1478 = (8'haa);
            end
        end
    end
  assign wire1479 = $unsigned($unsigned({$unsigned($signed(wire1435)),
                        $signed($signed(reg1440))}));
  assign wire1480 = $signed({(~^reg1460[(4'h8):(3'h6)]),
                        ($signed(wire1434) ?
                            ((reg1456 ?
                                reg1476 : reg1448) >>> (~|reg1457)) : (+(-(8'ha1))))});
  always
    @(posedge clk) begin
      reg1481 = reg1441;
      reg1482 = reg1450;
    end
  always
    @(posedge clk) begin
      reg1483 = ($unsigned((~&reg1448)) ?
          wire1433[(2'h3):(2'h2)] : $signed(reg1437));
      if ((~($signed({reg1437[(4'h8):(2'h3)]}) ?
          (^~reg1445[(4'h9):(3'h4)]) : (wire1464[(5'h13):(5'h12)] && (reg1460[(3'h4):(3'h4)] > $unsigned(reg1440))))))
        begin
          for (forvar1484 = (1'h0); (forvar1484 < (1'h0)); forvar1484 = (forvar1484 + (1'h1)))
            begin
              reg1485 <= {{wire1465}, wire1436};
              reg1486 <= (reg1440 <= {(^~$unsigned((wire1464 ?
                      reg1450 : wire1435))),
                  $unsigned(($unsigned(reg1450) ? (!(8'hb5)) : wire1479))});
            end
          reg1487 = (+(~^wire1464[(5'h10):(1'h1)]));
        end
      else
        begin
          reg1484 = (~|wire1436);
          if ((|$signed($signed((reg1476[(3'h4):(2'h2)] ?
              {(8'ha0)} : (wire1434 ? reg1437 : reg1485))))))
            begin
              reg1487 = ({$unsigned(reg1475), wire1464[(4'he):(1'h1)]} ?
                  $signed((reg1441[(4'ha):(2'h2)] - $unsigned(reg1450))) : wire1436);
              reg1488 = (reg1440 ?
                  wire1465[(4'ha):(2'h3)] : $signed(((8'hbb) < ($unsigned(wire1434) < (wire1465 + reg1442)))));
              reg1489 = reg1460[(1'h1):(1'h1)];
              reg1490 <= $signed($unsigned(({$unsigned(reg1457), (-reg1483)} ?
                  $unsigned(wire1434[(4'hb):(4'ha)]) : {(wire1479 > forvar1484),
                      (reg1475 * reg1484)})));
            end
          else
            begin
              reg1485 <= reg1456;
              reg1487 = ((reg1485[(4'hf):(1'h1)] ?
                      (~^(reg1488[(1'h0):(1'h0)] ?
                          $unsigned(reg1457) : reg1476[(4'h9):(3'h6)])) : (forvar1484[(1'h1):(1'h0)] <= $signed(wire1464))) ?
                  (8'hbe) : {(~&(^reg1487[(4'ha):(4'h8)])),
                      reg1439[(4'he):(2'h3)]});
              reg1490 <= wire1435;
            end
          if (reg1450[(4'ha):(1'h1)])
            begin
              reg1491 = reg1475;
              reg1492 = $signed((7'h44));
              reg1493 <= (($signed(((~^wire1436) ?
                      $signed(reg1438) : (reg1450 && reg1488))) ~^ (reg1483 == ((reg1460 > (7'h41)) ?
                      reg1458 : (reg1490 ? reg1487 : wire1434)))) ?
                  $unsigned($signed(reg1488[(4'hf):(4'h9)])) : $signed($signed(((reg1487 == reg1460) ?
                      reg1437[(5'h13):(1'h1)] : {wire1479}))));
            end
          else
            begin
              reg1491 = ($signed(reg1489[(4'h8):(1'h0)]) | reg1443);
            end
        end
    end
  always
    @(posedge clk) begin
      reg1494 <= $unsigned((|((|{(8'hb1)}) ?
          reg1457[(2'h3):(1'h0)] : (~^$unsigned(reg1493)))));
      if (reg1457[(2'h2):(1'h1)])
        begin
          reg1495 <= reg1486;
          reg1496 <= (reg1457[(3'h4):(1'h1)] >>> ($unsigned(reg1438[(2'h2):(2'h2)]) ?
              reg1486[(3'h7):(1'h1)] : $signed(reg1495)));
        end
      else
        begin
          reg1495 <= (reg1443[(1'h0):(1'h0)] == (wire1464[(1'h1):(1'h1)] ?
              $unsigned((7'h48)) : $unsigned({reg1443[(4'ha):(4'h9)]})));
          reg1497 = ($unsigned($signed($signed((reg1448 >= (8'hbb))))) ?
              (|reg1495) : $unsigned(wire1435));
          if (reg1496)
            begin
              reg1498 <= $signed(($unsigned({$signed(reg1458)}) ~^ reg1485));
              reg1499 = ((8'hbb) & (~^($signed($unsigned((7'h47))) ?
                  reg1450[(2'h2):(1'h0)] : ($unsigned(reg1443) ^ reg1476[(5'h10):(4'hc)]))));
              reg1500 = $signed({$unsigned($unsigned((wire1464 & wire1465))),
                  $unsigned((reg1439[(5'h11):(4'hc)] <= (wire1464 ?
                      wire1433 : wire1434)))});
            end
          else
            begin
              reg1499 = $unsigned((&(^~$signed($unsigned((7'h47))))));
              reg1500 = ($signed($signed($unsigned((8'hba)))) ?
                  reg1475 : ($unsigned((reg1442[(1'h0):(1'h0)] == $signed(reg1499))) ?
                      reg1458[(4'ha):(2'h2)] : (reg1485 <= ($signed(wire1435) <= reg1490[(1'h1):(1'h1)]))));
              reg1501 <= reg1445;
              reg1502 <= (^~(reg1475 ? reg1476 : reg1450[(4'hb):(2'h2)]));
              reg1503 = reg1500[(4'hb):(1'h0)];
            end
          for (forvar1504 = (1'h0); (forvar1504 < (1'h0)); forvar1504 = (forvar1504 + (1'h1)))
            begin
              reg1505 = (($unsigned(((reg1440 <<< reg1499) ?
                      $unsigned(reg1440) : reg1495[(3'h5):(2'h2)])) <= ($signed(forvar1504) - $unsigned((!(8'hac))))) ?
                  $signed($unsigned($signed((forvar1504 ?
                      reg1499 : (8'haf))))) : (8'hb6));
            end
        end
      if ($signed(reg1498))
        begin
          reg1506 <= (^~$unsigned(reg1502[(3'h4):(1'h0)]));
          if ({$signed((|reg1495))})
            begin
              reg1507 <= ($unsigned((({reg1457} ?
                  $unsigned(reg1502) : ((8'hb7) ?
                      (8'ha2) : reg1499)) ^ ({(8'h9c), wire1465} ?
                  {wire1464} : wire1464[(1'h1):(1'h0)]))) | (8'hb7));
              reg1508 <= $signed(($signed(reg1498[(4'he):(1'h1)]) == $unsigned(reg1486)));
              reg1509 = (^~reg1486[(4'ha):(2'h3)]);
              reg1510 <= (reg1507 < ((7'h45) >>> $signed((^(wire1435 <= reg1501)))));
            end
          else
            begin
              reg1507 <= $unsigned((~|reg1507));
              reg1509 = {reg1442, $unsigned($signed(reg1460))};
            end
        end
      else
        begin
          if ((reg1443[(1'h1):(1'h0)] <= ($unsigned(reg1450[(2'h3):(1'h0)]) ?
              {$signed($unsigned((8'hb6)))} : (&$unsigned((&reg1494))))))
            begin
              reg1509 = (8'hb6);
              reg1511 = $signed(((|$unsigned(reg1439)) ?
                  (!((reg1505 ?
                      wire1436 : wire1453) < reg1499)) : $unsigned($unsigned((reg1497 && reg1448)))));
              reg1512 = reg1476[(2'h2):(1'h0)];
              reg1513 <= $signed((8'ha9));
              reg1514 <= $signed(((|($unsigned(reg1497) | $unsigned(reg1458))) ?
                  (reg1494 == ((8'ha5) >= (~reg1476))) : reg1508[(1'h1):(1'h1)]));
            end
          else
            begin
              reg1506 <= $unsigned(($unsigned($unsigned((reg1458 ?
                      (8'ha7) : reg1502))) ?
                  reg1501 : $signed(wire1479[(3'h7):(3'h7)])));
            end
          for (forvar1515 = (1'h0); (forvar1515 < (1'h1)); forvar1515 = (forvar1515 + (1'h1)))
            begin
              reg1516 = ($signed($signed(reg1505)) <= wire1435[(4'h8):(3'h5)]);
              reg1517 = $signed((^{($signed(reg1448) + (reg1440 ?
                      reg1509 : reg1494)),
                  $signed((forvar1504 ? (8'hbb) : reg1500))}));
            end
          for (forvar1518 = (1'h0); (forvar1518 < (2'h3)); forvar1518 = (forvar1518 + (1'h1)))
            begin
              reg1519 <= ((!((~(|wire1479)) ?
                  ({reg1511} && (8'had)) : ((reg1512 ? (7'h41) : reg1476) ?
                      (reg1498 || reg1507) : $signed((8'ha6))))) ^ (reg1440 ?
                  $signed({(reg1437 - (8'hbf))}) : reg1458[(1'h0):(1'h0)]));
              reg1520 = (-$signed($unsigned(((&(7'h4a)) && (reg1494 ?
                  reg1442 : reg1512)))));
            end
        end
    end
  assign wire1521 = $signed(($unsigned($unsigned(reg1457)) << {$signed((reg1438 ?
                            reg1501 : reg1485))}));
  assign wire1522 = (+($signed((((8'h9d) ^~ (8'hb5)) ^ $signed(wire1435))) <= reg1485[(5'h10):(3'h7)]));
  assign wire1523 = ((~|$unsigned($unsigned((reg1485 >= reg1502)))) <<< $unsigned(reg1448));
  always
    @(posedge clk) begin
      reg1524 <= (reg1506[(5'h10):(4'he)] <= (-reg1442[(4'ha):(2'h2)]));
      if (((reg1514[(4'hc):(4'hc)] << (~$unsigned(reg1485))) ?
          (((~^wire1522) == ((7'h4a) ?
              (+reg1510) : (reg1508 << (7'h42)))) > (($unsigned(reg1495) ?
                  reg1458 : (wire1522 ? reg1475 : (8'hbc))) ?
              wire1521 : reg1445[(3'h5):(2'h2)])) : reg1524[(4'ha):(3'h7)]))
        begin
          for (forvar1525 = (1'h0); (forvar1525 < (3'h4)); forvar1525 = (forvar1525 + (1'h1)))
            begin
              reg1526 <= ((($unsigned((8'hb2)) + {(~|reg1486)}) ?
                  $unsigned($unsigned(reg1475)) : $signed($unsigned((+reg1442)))) <<< ($signed(reg1457) ~^ (reg1502[(3'h7):(2'h3)] ?
                  (reg1460[(3'h7):(2'h2)] != (!wire1465)) : (reg1514[(4'ha):(4'h8)] ^~ wire1522))));
              reg1527 <= $signed($signed(reg1437));
              reg1528 <= (reg1524 >> reg1445);
            end
          for (forvar1529 = (1'h0); (forvar1529 < (3'h4)); forvar1529 = (forvar1529 + (1'h1)))
            begin
              reg1530 <= reg1498;
              reg1531 = $signed($unsigned(wire1521));
            end
          reg1532 <= (&(+(~|$unsigned((|(8'haf))))));
          reg1533 <= {($unsigned((reg1493[(3'h6):(3'h6)] & reg1507[(1'h0):(1'h0)])) ?
                  $unsigned((reg1514[(3'h5):(3'h5)] ?
                      ((7'h4a) < (7'h42)) : reg1457[(1'h0):(1'h0)])) : (~$unsigned(reg1441))),
              (8'h9c)};
        end
      else
        begin
          for (forvar1525 = (1'h0); (forvar1525 < (2'h2)); forvar1525 = (forvar1525 + (1'h1)))
            begin
              reg1529 = (8'hb4);
            end
          for (forvar1530 = (1'h0); (forvar1530 < (2'h3)); forvar1530 = (forvar1530 + (1'h1)))
            begin
              reg1532 <= (~$signed(((&(reg1442 ?
                  forvar1530 : reg1513)) == $unsigned(reg1493[(1'h0):(1'h0)]))));
              reg1533 <= (8'ha8);
              reg1534 = ($unsigned(reg1508) != reg1513);
              reg1535 <= ($unsigned({reg1527,
                  forvar1525[(3'h6):(3'h6)]}) >>> $signed($unsigned({reg1527})));
            end
          reg1536 = reg1506[(2'h3):(1'h1)];
          for (forvar1537 = (1'h0); (forvar1537 < (2'h3)); forvar1537 = (forvar1537 + (1'h1)))
            begin
              reg1538 <= reg1533;
              reg1539 = ($signed((-reg1528[(2'h2):(1'h0)])) != $signed(reg1535[(4'ha):(3'h4)]));
              reg1540 = wire1434[(1'h1):(1'h0)];
              reg1541 <= (reg1513 ^~ (((|reg1443) ? reg1438 : forvar1529) ?
                  $unsigned((+(reg1538 ?
                      reg1494 : reg1440))) : $unsigned((^reg1506[(5'h13):(4'hb)]))));
              reg1542 <= reg1531;
            end
          reg1543 = (~(~&{(~wire1522), wire1433}));
        end
      if ((reg1456[(4'h9):(3'h7)] ?
          ($signed((+{reg1514, (8'h9f)})) ?
              {reg1457[(1'h0):(1'h0)],
                  (~&$signed(reg1539))} : (($signed(wire1464) <= (8'h9f)) + {$unsigned(wire1453)})) : $signed(wire1521)))
        begin
          if ($unsigned(reg1441))
            begin
              reg1544 = $signed(reg1486[(3'h7):(2'h2)]);
              reg1545 <= (reg1540[(1'h0):(1'h0)] ?
                  reg1457 : $signed($unsigned($signed((reg1458 ?
                      reg1542 : reg1510)))));
            end
          else
            begin
              reg1544 = (8'ha1);
              reg1546 = $signed($signed(reg1527[(3'h5):(1'h0)]));
              reg1547 <= (+reg1532[(4'h8):(1'h0)]);
            end
          if (reg1448)
            begin
              reg1548 <= reg1530;
              reg1549 <= {($unsigned((&(reg1524 ~^ reg1538))) ?
                      ((~&(wire1464 ?
                          forvar1530 : reg1439)) || $signed($signed(forvar1525))) : (($signed(forvar1537) >>> (reg1490 ?
                          (8'hae) : wire1480)) >= reg1486)),
                  (({(8'hbf),
                          (reg1495 >> (8'had))} >> (^reg1445[(5'h10):(3'h7)])) ?
                      $signed($unsigned($unsigned((8'hac)))) : reg1475)};
            end
          else
            begin
              reg1548 <= $unsigned(wire1433[(3'h4):(2'h3)]);
              reg1549 <= reg1439;
              reg1550 = $unsigned((reg1445[(5'h11):(3'h7)] - reg1529));
              reg1551 <= $signed(((7'h42) > $unsigned(({reg1460,
                  reg1545} >= reg1508))));
            end
          reg1552 = (($unsigned(wire1464) ?
              wire1435[(4'he):(2'h3)] : {(+reg1529)}) <<< ({($signed(reg1524) && {(8'hbf)})} ?
              (~&wire1435[(3'h6):(2'h2)]) : $signed(((reg1493 ?
                      wire1522 : wire1436) ?
                  reg1549[(4'ha):(4'h8)] : {reg1535, reg1494}))));
          for (forvar1553 = (1'h0); (forvar1553 < (1'h0)); forvar1553 = (forvar1553 + (1'h1)))
            begin
              reg1554 <= ((+(+reg1508)) ?
                  reg1490 : (&((8'ha9) <= ($unsigned(wire1453) ?
                      (reg1527 ? (8'h9f) : reg1543) : (~reg1476)))));
              reg1555 = (7'h44);
              reg1556 <= $unsigned(wire1465);
            end
          for (forvar1557 = (1'h0); (forvar1557 < (1'h0)); forvar1557 = (forvar1557 + (1'h1)))
            begin
              reg1558 <= ($unsigned($unsigned(((-reg1437) ?
                      (reg1445 ?
                          (7'h47) : (8'hbd)) : forvar1529[(2'h3):(1'h0)]))) ?
                  {{$signed((wire1434 ? wire1465 : reg1439)),
                          (reg1550[(2'h3):(1'h0)] & $signed(wire1435))}} : reg1437[(1'h0):(1'h0)]);
              reg1559 = ((-reg1501) ?
                  $unsigned(({reg1556[(2'h3):(1'h0)]} ?
                      (reg1457 >>> (forvar1529 ?
                          reg1526 : reg1538)) : reg1547[(3'h5):(2'h2)])) : reg1495[(4'hd):(4'hd)]);
              reg1560 = $signed($signed({(reg1442 >>> (reg1510 ?
                      reg1485 : reg1490))}));
            end
        end
      else
        begin
          reg1545 <= (reg1546[(4'hc):(3'h7)] ?
              reg1513[(1'h0):(1'h0)] : $unsigned(reg1441));
          for (forvar1546 = (1'h0); (forvar1546 < (2'h2)); forvar1546 = (forvar1546 + (1'h1)))
            begin
              reg1547 <= ((reg1514 ?
                      {forvar1525,
                          ($signed(forvar1553) <= (reg1476 + reg1549))} : (((reg1543 ^ reg1548) - (~^reg1441)) ?
                          $signed((-(8'hb0))) : reg1443)) ?
                  reg1448[(2'h3):(1'h0)] : ({reg1445,
                      ($unsigned(reg1438) ?
                          (wire1479 && reg1555) : (-reg1547))} ^~ {reg1529[(2'h3):(2'h3)]}));
              reg1548 <= reg1450;
              reg1549 <= (~^($unsigned((!$unsigned(reg1546))) ?
                  {$signed(reg1559),
                      ({reg1507, (8'hb5)} || reg1555)} : reg1450));
              reg1550 = ((reg1458 ?
                      ({(reg1493 ? reg1443 : reg1552), reg1528} ?
                          {(reg1544 == wire1433),
                              (reg1547 > forvar1525)} : $unsigned((reg1439 & reg1555))) : $unsigned($unsigned({reg1549}))) ?
                  reg1554[(2'h2):(2'h2)] : reg1535);
            end
          for (forvar1551 = (1'h0); (forvar1551 < (2'h2)); forvar1551 = (forvar1551 + (1'h1)))
            begin
              reg1553 <= {$signed((((reg1545 ?
                          reg1460 : (7'h44)) && ((7'h49) || reg1547)) ?
                      {(&reg1524)} : reg1545)),
                  (({(reg1552 ?
                          reg1476 : (8'ha2))} - $signed((reg1548 > wire1453))) != (!($unsigned(reg1458) ?
                      $signed(wire1480) : reg1531[(4'hc):(4'h8)])))};
            end
          reg1555 = wire1435[(3'h5):(2'h2)];
          for (forvar1556 = (1'h0); (forvar1556 < (1'h1)); forvar1556 = (forvar1556 + (1'h1)))
            begin
              reg1557 <= (^reg1508);
              reg1559 = $signed({$signed(($unsigned((8'hb6)) + $signed(reg1460)))});
              reg1561 <= reg1440[(2'h2):(1'h0)];
            end
        end
    end
  always
    @(posedge clk) begin
      reg1562 = reg1445;
    end
  assign wire1563 = ((reg1545[(4'he):(3'h5)] ?
                        wire1523 : (((-reg1493) & reg1442[(3'h7):(1'h0)]) & (8'ha6))) != reg1485[(5'h10):(3'h4)]);
  assign wire1564 = reg1475;
  always
    @(posedge clk) begin
      reg1565 = $unsigned(($signed(({reg1524, reg1502} <<< $signed((8'hb0)))) ?
          $unsigned({reg1524[(2'h2):(1'h0)], (8'haa)}) : reg1502));
      if ((reg1496 == $signed({reg1438})))
        begin
          if (wire1563[(4'h8):(3'h4)])
            begin
              reg1566 = ({(~(|(reg1490 ?
                      (8'hb4) : reg1526)))} > $signed(({$signed((8'ha6))} ?
                  $unsigned(reg1445[(4'hc):(1'h0)]) : {reg1533,
                      wire1563[(1'h1):(1'h1)]})));
              reg1567 <= reg1501;
              reg1568 = ((((&(-reg1514)) ?
                          reg1445 : $signed((reg1437 ? reg1437 : reg1501))) ?
                      (((&wire1523) || (^~reg1526)) ?
                          $unsigned(reg1549) : (~|(reg1439 ?
                              (8'hac) : reg1526))) : {(^~reg1557),
                          (!reg1519)}) ?
                  (~&(|reg1486)) : $signed($signed($signed((~&wire1563)))));
            end
          else
            begin
              reg1566 = (|(|reg1498));
              reg1567 <= reg1440;
              reg1568 = (wire1434[(2'h2):(2'h2)] ?
                  reg1551 : {(($unsigned(reg1440) << reg1553) ?
                          reg1475[(1'h1):(1'h0)] : reg1456[(1'h1):(1'h1)]),
                      reg1524[(1'h0):(1'h0)]});
            end
          if ($signed(($unsigned(reg1456) ?
              (~|$signed($signed(reg1441))) : $signed(((reg1508 >= reg1530) ?
                  reg1438[(2'h2):(1'h0)] : reg1567)))))
            begin
              reg1569 = (~&$signed($signed(($unsigned(wire1479) ^~ (reg1545 ?
                  reg1510 : reg1528)))));
              reg1570 = (8'hbb);
              reg1571 = $unsigned((!reg1554[(4'hd):(3'h6)]));
              reg1572 = $signed((wire1435[(4'ha):(3'h7)] < $signed(wire1480[(2'h3):(1'h0)])));
              reg1573 = (~&(^$unsigned((7'h45))));
            end
          else
            begin
              reg1574 <= $unsigned(({(-$unsigned(reg1551))} == reg1573));
              reg1575 = $signed($unsigned(((reg1441[(4'he):(4'ha)] >>> (reg1442 ?
                      (7'h48) : (8'hae))) ?
                  $signed((^reg1441)) : reg1566)));
              reg1576 = {($signed($signed(reg1565[(3'h7):(3'h5)])) ?
                      ($unsigned(reg1542) ?
                          reg1508[(1'h1):(1'h1)] : reg1548) : $unsigned(((reg1514 <= reg1507) != reg1569)))};
              reg1577 <= {reg1572[(4'hb):(4'ha)]};
            end
        end
      else
        begin
          reg1566 = $unsigned(reg1577[(4'ha):(4'h9)]);
          if ($signed(((+reg1524[(4'hd):(2'h3)]) | reg1494[(1'h0):(1'h0)])))
            begin
              reg1568 = ((^~reg1561[(3'h6):(2'h3)]) ~^ ((+(~^reg1514[(4'h9):(3'h5)])) ?
                  (|$signed((~^reg1519))) : reg1577));
            end
          else
            begin
              reg1567 <= (|reg1567[(3'h7):(2'h3)]);
            end
          reg1574 <= ($signed((7'h47)) ?
              ($unsigned((((8'ha4) & reg1510) >> $unsigned(reg1567))) && (reg1571 && reg1569)) : ((((!reg1498) || wire1564[(4'h8):(3'h4)]) ?
                      $unsigned((^~wire1564)) : reg1441) ?
                  reg1441[(3'h5):(1'h1)] : (($signed(reg1561) ?
                      $unsigned(reg1498) : {reg1445,
                          reg1494}) - ((reg1549 >>> reg1486) <<< (|(7'h48))))));
        end
      reg1578 <= (!reg1568[(4'h8):(3'h4)]);
      reg1579 <= (&{(~&(-reg1448[(2'h2):(1'h0)])), wire1479[(4'hb):(3'h4)]});
    end
  always
    @(posedge clk) begin
      reg1580 <= ($signed((((wire1564 ?
                  reg1442 : reg1476) && (reg1549 >> reg1440)) ?
              ($signed((8'hba)) ?
                  $signed(reg1443) : wire1523) : $unsigned({(8'hac),
                  reg1530}))) ?
          wire1464 : wire1521);
      for (forvar1581 = (1'h0); (forvar1581 < (2'h2)); forvar1581 = (forvar1581 + (1'h1)))
        begin
          if ($signed($signed(($unsigned(reg1556[(1'h0):(1'h0)]) ?
              reg1556[(3'h7):(2'h2)] : $unsigned((&reg1450))))))
            begin
              reg1582 = $signed($signed(($unsigned((reg1526 ~^ reg1578)) > (~^(^reg1542)))));
              reg1583 = $unsigned((~(|($unsigned(reg1578) ?
                  $signed((7'h48)) : $unsigned(reg1458)))));
              reg1584 = (!$unsigned((~(-(reg1442 & reg1579)))));
              reg1585 = (^~reg1439[(4'he):(3'h5)]);
            end
          else
            begin
              reg1582 = reg1507;
            end
          reg1586 = (((^$unsigned($unsigned(wire1522))) ?
              (~$signed(reg1475[(1'h0):(1'h0)])) : (|({wire1564, reg1495} ?
                  reg1443 : reg1548))) || reg1490);
          for (forvar1587 = (1'h0); (forvar1587 < (2'h2)); forvar1587 = (forvar1587 + (1'h1)))
            begin
              reg1588 <= reg1456;
              reg1589 = $unsigned((+(!((-reg1526) ?
                  (reg1485 ? reg1486 : reg1498) : (reg1501 <<< forvar1587)))));
              reg1590 = (|(reg1589 >= reg1586[(3'h4):(2'h3)]));
              reg1591 = reg1557;
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1142  (y, clk, wire1147, wire1146, wire1145, wire1144, wire1143);
  output wire [(32'h9e1):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire1147;
  input wire [(4'hd):(1'h0)] wire1146;
  input wire signed [(4'he):(1'h0)] wire1145;
  input wire signed [(4'ha):(1'h0)] wire1144;
  input wire signed [(5'h16):(1'h0)] wire1143;
  wire signed [(5'h11):(1'h0)] wire1266;
  wire signed [(2'h3):(1'h0)] wire1265;
  wire signed [(5'h16):(1'h0)] wire1264;
  wire [(4'hf):(1'h0)] wire1215;
  wire [(3'h4):(1'h0)] wire1214;
  wire [(5'h16):(1'h0)] wire1207;
  wire signed [(4'hd):(1'h0)] wire1206;
  wire signed [(4'ha):(1'h0)] wire1172;
  wire [(5'h16):(1'h0)] wire1171;
  wire signed [(3'h6):(1'h0)] wire1148;
  reg [(5'h12):(1'h0)] reg1333 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1332 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1331 = (1'h0);
  reg [(5'h17):(1'h0)] reg1325 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1321 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1314 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1309 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1305 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1304 = (1'h0);
  reg [(4'ha):(1'h0)] reg1301 = (1'h0);
  reg [(4'h8):(1'h0)] reg1300 = (1'h0);
  reg [(5'h14):(1'h0)] reg1299 = (1'h0);
  reg [(3'h4):(1'h0)] reg1297 = (1'h0);
  reg [(5'h16):(1'h0)] reg1295 = (1'h0);
  reg [(4'hd):(1'h0)] reg1293 = (1'h0);
  reg [(2'h3):(1'h0)] reg1291 = (1'h0);
  reg [(3'h6):(1'h0)] reg1285 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1284 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1281 = (1'h0);
  reg [(4'h9):(1'h0)] reg1280 = (1'h0);
  reg [(5'h15):(1'h0)] reg1278 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1275 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1274 = (1'h0);
  reg [(5'h13):(1'h0)] reg1269 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1259 = (1'h0);
  reg [(3'h6):(1'h0)] reg1257 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1256 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1253 = (1'h0);
  reg [(5'h18):(1'h0)] reg1250 = (1'h0);
  reg [(4'hc):(1'h0)] reg1249 = (1'h0);
  reg [(3'h6):(1'h0)] reg1248 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1237 = (1'h0);
  reg [(4'he):(1'h0)] reg1236 = (1'h0);
  reg [(4'hd):(1'h0)] reg1234 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1229 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1228 = (1'h0);
  reg [(5'h10):(1'h0)] reg1222 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1225 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1223 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1220 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1218 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1217 = (1'h0);
  reg [(5'h14):(1'h0)] reg1216 = (1'h0);
  reg [(5'h17):(1'h0)] reg1211 = (1'h0);
  reg [(4'h8):(1'h0)] reg1209 = (1'h0);
  reg [(4'hd):(1'h0)] reg1208 = (1'h0);
  reg [(5'h16):(1'h0)] reg1205 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1203 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1200 = (1'h0);
  reg [(5'h18):(1'h0)] reg1199 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1198 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1195 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1194 = (1'h0);
  reg [(4'hd):(1'h0)] reg1191 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1190 = (1'h0);
  reg [(5'h10):(1'h0)] reg1188 = (1'h0);
  reg [(5'h16):(1'h0)] reg1187 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1186 = (1'h0);
  reg [(5'h10):(1'h0)] reg1185 = (1'h0);
  reg [(5'h14):(1'h0)] reg1175 = (1'h0);
  reg [(5'h17):(1'h0)] reg1184 = (1'h0);
  reg [(4'h8):(1'h0)] reg1183 = (1'h0);
  reg [(5'h16):(1'h0)] reg1181 = (1'h0);
  reg [(4'hd):(1'h0)] reg1179 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1177 = (1'h0);
  reg [(5'h18):(1'h0)] reg1173 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1168 = (1'h0);
  reg [(2'h3):(1'h0)] reg1164 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1160 = (1'h0);
  reg [(5'h17):(1'h0)] reg1159 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1158 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1157 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1153 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1151 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1149 = (1'h0);
  reg [(3'h4):(1'h0)] reg1334 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1330 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1329 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1328 = (1'h0);
  reg [(2'h2):(1'h0)] reg1327 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1326 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1324 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1323 = (1'h0);
  reg [(5'h12):(1'h0)] reg1322 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1320 = (1'h0);
  reg [(3'h6):(1'h0)] reg1319 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1318 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1317 = (1'h0);
  reg [(5'h15):(1'h0)] reg1316 = (1'h0);
  reg [(4'h8):(1'h0)] reg1315 = (1'h0);
  reg [(4'hd):(1'h0)] reg1313 = (1'h0);
  reg [(5'h14):(1'h0)] reg1312 = (1'h0);
  reg [(3'h5):(1'h0)] reg1311 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1310 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1308 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1307 = (1'h0);
  reg [(5'h12):(1'h0)] reg1306 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1303 = (1'h0);
  reg [(4'h8):(1'h0)] reg1302 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1298 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1296 = (1'h0);
  reg [(4'h9):(1'h0)] reg1294 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1292 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1290 = (1'h0);
  reg [(4'hf):(1'h0)] reg1289 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1288 = (1'h0);
  reg [(3'h4):(1'h0)] reg1287 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1286 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1283 = (1'h0);
  reg [(5'h10):(1'h0)] reg1282 = (1'h0);
  reg [(5'h14):(1'h0)] reg1279 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1277 = (1'h0);
  reg [(4'ha):(1'h0)] reg1276 = (1'h0);
  reg [(5'h14):(1'h0)] reg1273 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1272 = (1'h0);
  reg [(2'h3):(1'h0)] reg1271 = (1'h0);
  reg [(4'ha):(1'h0)] reg1270 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1268 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1267 = (1'h0);
  reg [(3'h5):(1'h0)] reg1263 = (1'h0);
  reg [(5'h18):(1'h0)] reg1262 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1261 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1260 = (1'h0);
  reg [(4'he):(1'h0)] reg1258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1255 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1252 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1255 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1254 = (1'h0);
  reg [(3'h6):(1'h0)] reg1252 = (1'h0);
  reg [(5'h12):(1'h0)] reg1251 = (1'h0);
  reg [(5'h10):(1'h0)] reg1247 = (1'h0);
  reg [(3'h5):(1'h0)] reg1246 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1245 = (1'h0);
  reg [(5'h13):(1'h0)] reg1244 = (1'h0);
  reg [(4'hf):(1'h0)] reg1243 = (1'h0);
  reg [(3'h5):(1'h0)] reg1242 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1241 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1240 = (1'h0);
  reg [(5'h13):(1'h0)] reg1239 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1238 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1235 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1233 = (1'h0);
  reg [(5'h10):(1'h0)] reg1232 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1231 = (1'h0);
  reg [(4'hc):(1'h0)] reg1230 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1227 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1226 = (1'h0);
  reg [(5'h12):(1'h0)] reg1224 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1222 = (1'h0);
  reg [(3'h7):(1'h0)] reg1221 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1219 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1213 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1212 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1210 = (1'h0);
  reg [(4'h8):(1'h0)] reg1204 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1202 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1201 = (1'h0);
  reg [(5'h16):(1'h0)] reg1197 = (1'h0);
  reg [(5'h14):(1'h0)] reg1196 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1193 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1192 = (1'h0);
  reg [(5'h17):(1'h0)] reg1189 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1182 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1180 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1178 = (1'h0);
  reg [(4'he):(1'h0)] reg1176 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1175 = (1'h0);
  reg [(4'hc):(1'h0)] reg1174 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1170 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1169 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1167 = (1'h0);
  reg [(4'hb):(1'h0)] reg1166 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1165 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1163 = (1'h0);
  reg [(4'hc):(1'h0)] reg1162 = (1'h0);
  reg [(5'h10):(1'h0)] reg1161 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1156 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1155 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1154 = (1'h0);
  reg [(4'h8):(1'h0)] reg1152 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1150 = (1'h0);
  assign y = {wire1266,
                 wire1265,
                 wire1264,
                 wire1215,
                 wire1214,
                 wire1207,
                 wire1206,
                 wire1172,
                 wire1171,
                 wire1148,
                 reg1333,
                 reg1332,
                 reg1331,
                 reg1325,
                 reg1321,
                 reg1314,
                 reg1309,
                 reg1305,
                 reg1304,
                 reg1301,
                 reg1300,
                 reg1299,
                 reg1297,
                 reg1295,
                 reg1293,
                 reg1291,
                 reg1285,
                 reg1284,
                 reg1281,
                 reg1280,
                 reg1278,
                 reg1275,
                 reg1274,
                 reg1269,
                 reg1259,
                 reg1257,
                 reg1256,
                 reg1253,
                 reg1250,
                 reg1249,
                 reg1248,
                 reg1237,
                 reg1236,
                 reg1234,
                 reg1229,
                 reg1228,
                 reg1222,
                 reg1225,
                 reg1223,
                 reg1220,
                 reg1218,
                 reg1217,
                 reg1216,
                 reg1211,
                 reg1209,
                 reg1208,
                 reg1205,
                 reg1203,
                 reg1200,
                 reg1199,
                 reg1198,
                 reg1195,
                 reg1194,
                 reg1191,
                 reg1190,
                 reg1188,
                 reg1187,
                 reg1186,
                 reg1185,
                 reg1175,
                 reg1184,
                 reg1183,
                 reg1181,
                 reg1179,
                 reg1177,
                 reg1173,
                 reg1168,
                 reg1164,
                 reg1160,
                 reg1159,
                 reg1158,
                 reg1157,
                 reg1153,
                 reg1151,
                 reg1149,
                 reg1334,
                 reg1330,
                 forvar1329,
                 reg1328,
                 reg1327,
                 forvar1326,
                 reg1324,
                 forvar1323,
                 reg1322,
                 reg1320,
                 reg1319,
                 forvar1318,
                 forvar1317,
                 reg1316,
                 reg1315,
                 reg1313,
                 reg1312,
                 reg1311,
                 reg1310,
                 forvar1308,
                 forvar1307,
                 reg1306,
                 forvar1303,
                 reg1302,
                 forvar1298,
                 reg1296,
                 reg1294,
                 forvar1292,
                 reg1290,
                 reg1289,
                 forvar1288,
                 reg1287,
                 reg1286,
                 reg1283,
                 reg1282,
                 reg1279,
                 reg1277,
                 reg1276,
                 reg1273,
                 reg1272,
                 reg1271,
                 reg1270,
                 forvar1268,
                 forvar1267,
                 reg1263,
                 reg1262,
                 reg1261,
                 forvar1260,
                 reg1258,
                 reg1255,
                 forvar1252,
                 forvar1255,
                 reg1254,
                 reg1252,
                 reg1251,
                 reg1247,
                 reg1246,
                 reg1245,
                 reg1244,
                 reg1243,
                 reg1242,
                 reg1241,
                 reg1240,
                 reg1239,
                 forvar1238,
                 forvar1235,
                 reg1233,
                 reg1232,
                 reg1231,
                 reg1230,
                 reg1227,
                 reg1226,
                 reg1224,
                 forvar1222,
                 reg1221,
                 reg1219,
                 reg1213,
                 reg1212,
                 reg1210,
                 reg1204,
                 reg1202,
                 reg1201,
                 reg1197,
                 reg1196,
                 reg1193,
                 forvar1192,
                 reg1189,
                 reg1182,
                 forvar1180,
                 reg1178,
                 reg1176,
                 forvar1175,
                 reg1174,
                 reg1170,
                 reg1169,
                 reg1167,
                 reg1166,
                 reg1165,
                 reg1163,
                 reg1162,
                 reg1161,
                 reg1156,
                 reg1155,
                 reg1154,
                 reg1152,
                 forvar1150,
                 (1'h0)};
  assign wire1148 = wire1145;
  always
    @(posedge clk) begin
      reg1149 <= $unsigned((($unsigned(wire1143[(5'h10):(5'h10)]) ?
              $unsigned(wire1146) : wire1143[(4'hc):(3'h4)]) ?
          (wire1144 ?
              ($signed(wire1143) & (|wire1144)) : $unsigned(wire1146)) : (wire1145[(4'hb):(4'hb)] < (wire1145 ^~ (7'h48)))));
      for (forvar1150 = (1'h0); (forvar1150 < (1'h1)); forvar1150 = (forvar1150 + (1'h1)))
        begin
          if (($signed(((|wire1144[(3'h7):(3'h5)]) ?
                  $signed((&(7'h42))) : (-$signed((7'h48))))) ?
              (&wire1147[(3'h6):(1'h1)]) : $unsigned((wire1146[(4'ha):(1'h1)] | wire1146[(4'hb):(4'hb)]))))
            begin
              reg1151 <= reg1149;
              reg1152 = wire1144;
              reg1153 <= reg1149[(4'ha):(3'h4)];
            end
          else
            begin
              reg1152 = reg1151;
              reg1154 = (8'had);
            end
          reg1155 = {wire1144[(1'h0):(1'h0)],
              $unsigned($unsigned($signed(reg1153[(1'h0):(1'h0)])))};
        end
      reg1156 = $unsigned((^~$unsigned($signed((reg1155 ?
          wire1144 : reg1152)))));
      if ($signed($unsigned(wire1146[(4'ha):(2'h2)])))
        begin
          reg1157 <= $signed((&((~^reg1153[(2'h3):(2'h2)]) ?
              $unsigned(reg1155) : wire1147)));
          reg1158 <= (reg1155[(2'h3):(1'h1)] ?
              ((({wire1145} ?
                  $unsigned(reg1149) : reg1152[(3'h6):(3'h4)]) & (~|(reg1153 <= reg1157))) != ((reg1154[(1'h1):(1'h1)] << (wire1145 + wire1145)) == ($unsigned(reg1156) ?
                  (|wire1148) : (reg1155 ?
                      reg1149 : reg1153)))) : ((reg1154 <<< {reg1151[(1'h1):(1'h1)],
                      wire1145}) ?
                  {(+wire1145[(3'h5):(3'h4)])} : {reg1151}));
          reg1159 <= wire1143;
          if (reg1158)
            begin
              reg1160 <= (((($unsigned(reg1154) << (reg1155 ?
                  reg1156 : forvar1150)) - $signed($unsigned(wire1144))) && (+{$signed((8'hac)),
                  (reg1159 <= wire1148)})) * $signed(reg1151));
              reg1161 = ((&$unsigned((reg1156[(5'h10):(4'hc)] ?
                      (wire1146 ^ reg1149) : $unsigned(reg1158)))) ?
                  $signed(reg1152) : (reg1151[(4'hf):(2'h2)] >> (+({wire1145} ?
                      $signed(wire1148) : $unsigned(reg1151)))));
              reg1162 = (8'haa);
              reg1163 = ((~^(~|forvar1150)) ^ ($signed(((|reg1153) ?
                      (~^wire1147) : (reg1155 >>> reg1161))) ?
                  (^~reg1154[(1'h1):(1'h1)]) : {{reg1152[(3'h7):(3'h7)],
                          (reg1159 ^~ wire1144)}}));
            end
          else
            begin
              reg1160 <= $signed({(reg1155 >= ({reg1155,
                      reg1163} == (8'hb4)))});
              reg1164 <= ($unsigned(reg1163) == ((reg1160 >> (7'h44)) >>> reg1161[(3'h7):(2'h2)]));
              reg1165 = (+$unsigned(((8'ha6) ? (^(^reg1161)) : wire1148)));
              reg1166 = {($signed($unsigned({reg1164, wire1145})) ?
                      (+reg1162) : $unsigned(wire1144))};
              reg1167 = reg1163;
            end
        end
      else
        begin
          if (((!$signed(wire1146[(3'h7):(3'h4)])) ? (8'h9c) : reg1158))
            begin
              reg1157 <= (|$signed(($signed(reg1161) ^~ ({reg1151} & (reg1154 ~^ (8'h9c))))));
              reg1158 <= (reg1163 ?
                  (^$unsigned(({reg1160, wire1148} ?
                      reg1166 : wire1148[(1'h1):(1'h1)]))) : ($signed(({reg1165} ?
                      $signed(reg1155) : (wire1146 ?
                          reg1149 : reg1165))) <= reg1154));
              reg1159 <= ((-((!reg1156) ?
                  reg1165 : ((|(8'hb9)) <= reg1161))) < (~&$unsigned((~^$unsigned((7'h40))))));
              reg1161 = forvar1150;
              reg1164 <= (+(+reg1160));
            end
          else
            begin
              reg1161 = $unsigned(((+$unsigned($unsigned(reg1160))) ?
                  forvar1150[(4'hf):(1'h0)] : ($signed(((8'ha1) - wire1144)) ?
                      (!(reg1166 ? reg1163 : reg1160)) : (~^(forvar1150 ?
                          wire1147 : (7'h46))))));
              reg1164 <= reg1152;
              reg1168 <= reg1166[(1'h1):(1'h1)];
            end
          reg1169 = {$signed((^reg1159))};
        end
      reg1170 = $signed($unsigned((reg1167 ?
          ((reg1154 ? reg1159 : reg1159) <<< (reg1165 ?
              reg1166 : reg1158)) : reg1162)));
    end
  assign wire1171 = wire1143[(5'h16):(2'h3)];
  assign wire1172 = $signed(({wire1147,
                        ($unsigned(wire1171) >> (wire1144 ?
                            reg1164 : reg1158))} * (7'h42)));
  always
    @(posedge clk) begin
      if ((wire1172[(3'h7):(3'h5)] ?
          {$signed($signed((reg1158 <<< reg1151)))} : {reg1149,
              $signed((reg1158[(2'h2):(2'h2)] ?
                  (~reg1164) : reg1159[(5'h12):(4'hb)]))}))
        begin
          reg1173 <= ($unsigned((!wire1171)) ?
              (((~|reg1149) ^~ reg1157[(4'ha):(4'h9)]) < $signed($unsigned({reg1168}))) : reg1158);
          reg1174 = $signed((8'hbf));
          for (forvar1175 = (1'h0); (forvar1175 < (3'h4)); forvar1175 = (forvar1175 + (1'h1)))
            begin
              reg1176 = (~&$signed($signed(reg1168)));
              reg1177 <= wire1172;
              reg1178 = $unsigned($signed(reg1149));
              reg1179 <= $signed(reg1157);
            end
          for (forvar1180 = (1'h0); (forvar1180 < (2'h2)); forvar1180 = (forvar1180 + (1'h1)))
            begin
              reg1181 <= (&$signed(((reg1173 ~^ (reg1174 ?
                      reg1168 : wire1148)) ?
                  $unsigned($signed(wire1144)) : $signed(reg1168))));
              reg1182 = ({$signed({(reg1164 ? wire1148 : reg1173)})} ?
                  $signed(reg1177[(4'h9):(4'h9)]) : $signed((!$signed(reg1149))));
              reg1183 <= $signed(($signed(reg1178[(4'he):(3'h6)]) <<< $unsigned(wire1145)));
              reg1184 <= (~^reg1174);
            end
        end
      else
        begin
          if (reg1183)
            begin
              reg1174 = $unsigned(({reg1157} ?
                  (~|$unsigned({reg1183})) : (((reg1179 ?
                          reg1158 : wire1172) | (|forvar1175)) ?
                      reg1160 : (wire1144 ? (7'h45) : (+reg1176)))));
            end
          else
            begin
              reg1174 = ((($signed(reg1159[(4'h9):(3'h6)]) ?
                      {$unsigned(reg1158),
                          (|reg1182)} : ((reg1160 <= reg1149) <= reg1158)) << (reg1164 & (8'haf))) ?
                  wire1171 : $unsigned((reg1157 ?
                      (~^forvar1180[(4'h9):(2'h3)]) : ($signed(wire1147) ?
                          (|(8'hbb)) : {wire1147}))));
            end
          reg1175 <= $signed({{(&(reg1160 ? reg1174 : reg1164))}});
        end
      if (forvar1175[(1'h1):(1'h0)])
        begin
          if (reg1164[(1'h0):(1'h0)])
            begin
              reg1185 <= $signed(reg1183);
              reg1186 <= (((({wire1147} ?
                      $signed(reg1177) : (^~reg1173)) && {(reg1177 ?
                          reg1176 : reg1157),
                      (reg1177 ?
                          (8'hb5) : reg1184)}) < reg1174[(3'h4):(1'h0)]) ?
                  wire1171[(4'he):(2'h2)] : (wire1144 ?
                      (((|(8'ha5)) | (wire1148 <= reg1185)) ?
                          reg1184 : (reg1183 < reg1178)) : $signed($unsigned((reg1151 ?
                          reg1178 : wire1146)))));
              reg1187 <= (7'h46);
              reg1188 <= (~&$signed(((~(reg1173 ?
                  wire1147 : reg1176)) == $unsigned(reg1168))));
            end
          else
            begin
              reg1189 = (forvar1175[(4'he):(3'h6)] == (^~$unsigned(reg1159[(1'h0):(1'h0)])));
            end
        end
      else
        begin
          if (($signed((((+(8'ha0)) + {reg1151}) | ((8'hb9) && {reg1175}))) < reg1178[(3'h5):(2'h2)]))
            begin
              reg1189 = ($unsigned({$unsigned((forvar1180 ?
                      wire1147 : wire1147)),
                  $unsigned(((8'hba) && reg1185))}) && ($unsigned(reg1184) ?
                  (|(~|(wire1148 <= reg1177))) : (~^((^wire1143) ?
                      $unsigned(reg1153) : $signed(wire1144)))));
              reg1190 <= (~^$signed(wire1171));
            end
          else
            begin
              reg1189 = $signed({($unsigned((reg1168 + reg1159)) ?
                      (8'hbb) : (-(reg1182 ? reg1187 : (7'h47))))});
            end
        end
      reg1191 <= $signed($signed($unsigned(($unsigned(reg1159) ?
          {wire1145} : $unsigned(wire1147)))));
      for (forvar1192 = (1'h0); (forvar1192 < (3'h4)); forvar1192 = (forvar1192 + (1'h1)))
        begin
          if ($unsigned($signed(reg1191)))
            begin
              reg1193 = (reg1164[(2'h3):(2'h3)] ?
                  ((((reg1178 <<< reg1177) <= {reg1191,
                          wire1145}) ^ {(reg1186 <<< wire1146)}) ?
                      $unsigned($unsigned(reg1184)) : reg1173[(4'hd):(1'h0)]) : (reg1149 ?
                      (~forvar1175) : ((~^(reg1157 + wire1143)) >>> {(reg1159 ?
                              reg1190 : (7'h4a)),
                          (+reg1190)})));
              reg1194 <= $unsigned((reg1191 ? forvar1180 : reg1182));
              reg1195 <= (-($unsigned($unsigned(reg1149[(5'h14):(4'h9)])) ?
                  (~{reg1188}) : (~^{(|reg1177)})));
            end
          else
            begin
              reg1194 <= ((|$signed((^~(7'h44)))) < $unsigned(($signed($signed(reg1195)) ?
                  (reg1191 ?
                      (reg1168 ?
                          reg1183 : wire1148) : wire1171[(5'h14):(3'h6)]) : $unsigned(((7'h4a) * reg1174)))));
              reg1196 = $unsigned($unsigned(reg1151[(4'hd):(4'h9)]));
            end
          reg1197 = ($signed(forvar1175[(4'h8):(3'h7)]) + wire1146);
          if (wire1171)
            begin
              reg1198 <= reg1186[(1'h0):(1'h0)];
              reg1199 <= reg1177;
              reg1200 <= wire1143[(5'h14):(1'h0)];
            end
          else
            begin
              reg1198 <= ((((~|$signed((8'ha1))) ?
                      (~&(-(8'hac))) : $unsigned(reg1173[(5'h13):(4'ha)])) > $signed($unsigned((reg1173 ?
                      (7'h42) : forvar1192)))) ?
                  reg1178[(4'h9):(3'h4)] : $signed(reg1149[(3'h5):(1'h0)]));
            end
          if (reg1174[(3'h7):(3'h5)])
            begin
              reg1201 = ($signed($unsigned((reg1188[(4'h9):(2'h2)] ?
                      ((7'h46) ^ forvar1192) : ((8'hb0) ?
                          reg1189 : wire1143)))) ?
                  (^$signed(reg1195[(5'h17):(4'ha)])) : (($unsigned((reg1198 ?
                          (8'had) : (7'h47))) <<< $signed(reg1159[(5'h10):(4'hf)])) ?
                      $unsigned(($unsigned(wire1146) ?
                          (wire1143 - forvar1192) : (wire1144 <<< reg1197))) : (7'h40)));
              reg1202 = {($unsigned({(reg1185 ? reg1195 : wire1172),
                      $unsigned((7'h40))}) - {reg1190[(1'h1):(1'h0)],
                      (reg1196[(1'h0):(1'h0)] <<< (reg1186 ?
                          wire1143 : reg1200))})};
            end
          else
            begin
              reg1203 <= {reg1186,
                  $unsigned((^~$unsigned((wire1143 <= reg1189))))};
            end
        end
      if ($unsigned(reg1191[(4'h8):(4'h8)]))
        begin
          reg1204 = {((^~$signed(((8'hb0) ? reg1173 : (8'hb4)))) ?
                  reg1198 : $signed({(+reg1184)})),
              {reg1198[(2'h2):(2'h2)],
                  $signed((|(reg1151 ? forvar1175 : reg1175)))}};
        end
      else
        begin
          reg1205 <= (reg1190 >= $signed($signed($signed(forvar1192))));
        end
    end
  assign wire1206 = (reg1160[(2'h2):(1'h0)] ?
                        $unsigned($signed(((wire1148 >>> wire1147) ?
                            reg1183[(3'h7):(1'h1)] : reg1157[(3'h4):(2'h2)]))) : {wire1145,
                            ((~^$unsigned(reg1173)) >> (&(!reg1173)))});
  assign wire1207 = $unsigned(reg1183);
  always
    @(posedge clk) begin
      reg1208 <= (reg1160[(3'h4):(3'h4)] ?
          $unsigned((reg1168[(2'h2):(2'h2)] | (+{reg1151,
              wire1145}))) : ({$signed({reg1153,
                  (8'ha0)})} <<< (($signed(reg1184) >> (+reg1190)) ?
              (^~{wire1172}) : (reg1185 ?
                  reg1185[(4'hc):(2'h3)] : $unsigned(reg1191)))));
      if ({$unsigned($unsigned((8'hbb)))})
        begin
          if (reg1173[(4'hb):(4'h9)])
            begin
              reg1209 <= (((!$unsigned((reg1173 ?
                  reg1195 : reg1179))) && (&$unsigned((reg1160 ?
                  wire1147 : wire1171)))) ^ wire1144[(3'h6):(3'h5)]);
              reg1210 = reg1190[(1'h1):(1'h0)];
              reg1211 <= $signed(reg1159);
              reg1212 = (reg1211 >>> {wire1147});
            end
          else
            begin
              reg1210 = $signed((reg1209[(2'h2):(1'h0)] >= $unsigned($signed(reg1153[(2'h2):(1'h0)]))));
              reg1211 <= (~|(reg1186[(3'h6):(3'h6)] ?
                  $signed(reg1190[(4'ha):(3'h5)]) : ((~^$unsigned(reg1157)) - reg1195[(5'h11):(3'h6)])));
              reg1212 = reg1181;
            end
          reg1213 = reg1159[(5'h17):(5'h14)];
        end
      else
        begin
          if ((({(~|((8'haf) ?
                      wire1206 : (8'hac)))} > ({wire1143[(1'h1):(1'h1)]} - $unsigned(reg1177[(3'h5):(1'h1)]))) ?
              {($signed($unsigned(reg1203)) ^ (^$unsigned((8'hb2)))),
                  ((^~reg1200) ?
                      reg1159 : ((+reg1160) ~^ {reg1158}))} : ({reg1153} ?
                  (~^reg1210[(3'h7):(2'h3)]) : {$signed((^(7'h45))),
                      $unsigned($signed(reg1194))})))
            begin
              reg1209 <= {(8'hbe),
                  $signed($unsigned($unsigned($signed(reg1190))))};
            end
          else
            begin
              reg1210 = reg1181;
              reg1211 <= $signed((reg1212[(3'h5):(1'h0)] > (($unsigned(reg1200) ?
                  ((8'hb5) ?
                      reg1210 : reg1164) : $signed(reg1186)) ^~ ((&wire1172) ?
                  (~&reg1181) : {reg1173}))));
            end
        end
    end
  assign wire1214 = wire1144[(3'h6):(1'h1)];
  assign wire1215 = $signed($signed(((8'hac) + {(~^wire1143)})));
  always
    @(posedge clk) begin
      if (reg1205[(5'h13):(3'h7)])
        begin
          reg1216 <= {(^~((|$signed(reg1175)) ?
                  {$unsigned(reg1211)} : $unsigned(reg1194))),
              (wire1147 ?
                  wire1206[(4'h9):(3'h4)] : $unsigned($signed({reg1151})))};
          if ($unsigned(wire1206[(3'h6):(2'h3)]))
            begin
              reg1217 <= $unsigned($unsigned((8'hb7)));
              reg1218 <= (reg1153[(3'h4):(1'h1)] ^~ $signed($signed($signed(reg1164[(2'h2):(2'h2)]))));
              reg1219 = (wire1146 ?
                  (^(!(reg1168 <<< (reg1211 ~^ reg1181)))) : wire1207[(1'h0):(1'h0)]);
              reg1220 <= $signed((((reg1168 ? $signed(reg1173) : reg1216) ?
                  reg1198[(2'h2):(1'h0)] : $unsigned((!(7'h46)))) << {({wire1146} ^ (wire1214 * reg1168))}));
              reg1221 = reg1198;
            end
          else
            begin
              reg1217 <= (reg1186 ?
                  {{reg1209, {(7'h40)}}} : (~&(~&$signed(reg1200))));
              reg1219 = reg1164[(1'h1):(1'h1)];
            end
          for (forvar1222 = (1'h0); (forvar1222 < (2'h2)); forvar1222 = (forvar1222 + (1'h1)))
            begin
              reg1223 <= $signed(reg1160);
              reg1224 = {(reg1195[(5'h16):(4'hb)] && (+{reg1164}))};
              reg1225 <= wire1147[(4'ha):(3'h7)];
              reg1226 = (((reg1175[(4'hd):(1'h0)] <= wire1171[(5'h16):(4'hd)]) ^~ reg1159[(4'hc):(4'h9)]) != reg1224);
            end
          reg1227 = reg1190[(2'h2):(1'h0)];
        end
      else
        begin
          reg1219 = ($signed((((~reg1177) >= reg1218) ~^ $unsigned($signed(wire1147)))) && (reg1200[(4'he):(4'ha)] ?
              (+(8'hac)) : {($unsigned(wire1206) ?
                      $signed(reg1221) : (reg1195 ? reg1220 : reg1203)),
                  ((reg1164 && wire1147) * wire1148)}));
          if (({{$signed($signed(reg1226))}} ?
              (reg1217[(2'h2):(1'h1)] ?
                  ($unsigned($unsigned(reg1160)) ?
                      (8'hbb) : $unsigned((reg1191 ?
                          reg1173 : wire1206))) : (^~((reg1151 - reg1188) ?
                      (^reg1187) : $unsigned(reg1217)))) : (reg1218[(3'h4):(1'h1)] ?
                  {wire1145} : reg1217)))
            begin
              reg1220 <= forvar1222;
              reg1222 <= reg1149;
              reg1223 <= (reg1225 + ($unsigned((((8'hbc) >= (8'hb4)) ?
                      (wire1146 << reg1223) : (~wire1215))) ?
                  reg1168[(4'he):(2'h3)] : $signed(reg1186[(1'h0):(1'h0)])));
            end
          else
            begin
              reg1221 = $signed({(~&(8'h9f)), (8'hb4)});
              reg1224 = reg1222;
              reg1225 <= (reg1185[(5'h10):(4'hb)] ?
                  (^{(wire1214[(1'h1):(1'h1)] ? {reg1158} : $signed((7'h47))),
                      ({reg1153, wire1206} ?
                          (reg1218 >>> wire1144) : reg1220[(2'h3):(2'h2)])}) : (~|$unsigned((^$signed(reg1158)))));
              reg1228 <= $signed((|reg1205));
            end
          if ($signed(reg1190))
            begin
              reg1229 <= ((((reg1186[(2'h2):(1'h0)] ?
                              $signed(reg1159) : reg1224[(3'h5):(1'h0)]) ?
                          ((wire1147 ? reg1217 : reg1223) ?
                              reg1168 : (|reg1199)) : $unsigned($signed(reg1168))) ?
                      reg1195 : $signed(({wire1172, reg1217} ?
                          $signed(reg1159) : $signed(reg1191)))) ?
                  reg1187[(3'h5):(1'h1)] : reg1187[(5'h12):(5'h10)]);
            end
          else
            begin
              reg1230 = wire1172[(3'h4):(1'h0)];
              reg1231 = reg1225[(1'h1):(1'h0)];
            end
          reg1232 = ((~&(-reg1153)) != reg1211);
        end
      reg1233 = $unsigned($unsigned(reg1177));
      reg1234 <= reg1232[(2'h3):(2'h3)];
    end
  always
    @(posedge clk) begin
      for (forvar1235 = (1'h0); (forvar1235 < (1'h0)); forvar1235 = (forvar1235 + (1'h1)))
        begin
          reg1236 <= wire1145;
          reg1237 <= reg1223;
        end
    end
  always
    @(posedge clk) begin
      for (forvar1238 = (1'h0); (forvar1238 < (2'h3)); forvar1238 = (forvar1238 + (1'h1)))
        begin
          reg1239 = (~&($unsigned($unsigned((wire1145 <<< reg1185))) ?
              reg1236[(1'h0):(1'h0)] : (&$unsigned((8'hb7)))));
          if (($unsigned($signed(reg1208)) ?
              (&(reg1218 <= {$signed(reg1239),
                  $signed(wire1207)})) : reg1177[(3'h7):(3'h7)]))
            begin
              reg1240 = (8'hb4);
              reg1241 = {$unsigned($unsigned($unsigned((reg1159 & reg1209)))),
                  ((&reg1236) || (~^((reg1153 ^~ wire1144) ?
                      (reg1157 ? reg1228 : wire1214) : {(7'h43), reg1209})))};
            end
          else
            begin
              reg1240 = (reg1217 ?
                  reg1240[(2'h3):(1'h1)] : reg1194[(2'h2):(1'h1)]);
              reg1241 = reg1186;
              reg1242 = reg1216[(2'h3):(1'h1)];
              reg1243 = ($signed(reg1183[(4'h8):(3'h6)]) ~^ (((reg1157 ?
                  (8'had) : (reg1236 ~^ reg1188)) - {(-reg1149)}) == wire1148));
              reg1244 = (!(!$signed((~&$signed((7'h48))))));
            end
        end
      reg1245 = (!(reg1173 <= $signed({(^~reg1151)})));
      if ((8'hb5))
        begin
          reg1246 = reg1199[(5'h18):(3'h4)];
          reg1247 = (!reg1195);
        end
      else
        begin
          reg1248 <= reg1203[(2'h3):(2'h2)];
        end
      if ($signed((reg1229[(1'h0):(1'h0)] ^ {$signed((7'h44))})))
        begin
          reg1249 <= reg1151;
          if (($unsigned(($unsigned((+reg1188)) ?
              wire1172 : $unsigned($signed((8'ha1))))) & $unsigned($signed({reg1243,
              (reg1191 * reg1177)}))))
            begin
              reg1250 <= $unsigned(reg1173[(5'h11):(3'h7)]);
              reg1251 = ((($unsigned((reg1187 + reg1236)) - (reg1190 ?
                      wire1144 : (reg1175 ? (8'ha9) : (7'h4a)))) ?
                  $signed(((~|reg1246) >>> (wire1148 != reg1228))) : $unsigned($signed(((8'haf) ^ reg1151)))) >> $signed(reg1246));
              reg1252 = $unsigned((^$signed(forvar1238)));
            end
          else
            begin
              reg1251 = reg1222;
              reg1253 <= wire1215;
            end
          reg1254 = ((|reg1240[(2'h3):(1'h0)]) ?
              $signed(((wire1207 > (reg1168 >= (8'ha6))) ?
                  reg1229[(3'h4):(2'h3)] : (((8'ha9) - wire1147) ?
                      (reg1190 ^ wire1147) : (8'ha6)))) : $signed((|$signed(reg1199[(4'h9):(4'h9)]))));
          for (forvar1255 = (1'h0); (forvar1255 < (1'h0)); forvar1255 = (forvar1255 + (1'h1)))
            begin
              reg1256 <= (($unsigned((8'ha2)) - ($signed(reg1205) ?
                  {(reg1225 ?
                          reg1200 : reg1246)} : ((reg1252 >>> (8'ha5)) | {wire1148,
                      wire1145}))) != (reg1149 ?
                  (reg1187 ?
                      $signed((8'ha7)) : (|reg1179)) : $unsigned((&$signed(forvar1238)))));
              reg1257 <= $signed(reg1234[(4'h8):(4'h8)]);
            end
        end
      else
        begin
          reg1251 = {(((~&$signed(reg1241)) ?
                  {(8'ha0),
                      $unsigned((8'hbd))} : reg1234) >>> (($signed(reg1239) + reg1241) ?
                  reg1199 : reg1228[(3'h4):(1'h1)]))};
          for (forvar1252 = (1'h0); (forvar1252 < (1'h1)); forvar1252 = (forvar1252 + (1'h1)))
            begin
              reg1253 <= ($signed((8'hbf)) ?
                  {(($signed(reg1203) ?
                          $signed(forvar1255) : $signed(reg1159)) ~^ $signed(reg1220[(1'h0):(1'h0)])),
                      $unsigned(((reg1220 * reg1211) ~^ $unsigned(reg1188)))} : $signed($unsigned($signed($unsigned((8'hb4))))));
              reg1254 = reg1157[(2'h3):(1'h1)];
              reg1255 = (forvar1255[(1'h1):(1'h0)] ?
                  ((^~((~reg1225) < $unsigned(reg1252))) ^ ({{reg1229}} != reg1168)) : wire1206);
              reg1258 = $signed(($signed((^(~&reg1157))) - reg1240[(1'h0):(1'h0)]));
            end
          reg1259 <= $signed(wire1144);
          for (forvar1260 = (1'h0); (forvar1260 < (2'h2)); forvar1260 = (forvar1260 + (1'h1)))
            begin
              reg1261 = wire1171[(4'h8):(1'h1)];
            end
          reg1262 = $unsigned((reg1239 != reg1244));
        end
    end
  always
    @(posedge clk) begin
      reg1263 = ((-$signed(reg1181)) ? reg1205[(3'h7):(1'h0)] : reg1218);
    end
  assign wire1264 = {{(reg1222[(4'h8):(2'h3)] ?
                                {(^(8'hbf))} : $signed((reg1188 > reg1208))),
                            (((!reg1200) ?
                                    (reg1203 + reg1217) : (reg1225 >> (8'ha6))) ?
                                ($unsigned(reg1149) ?
                                    $signed(reg1218) : $signed(wire1172)) : $signed((reg1234 <= reg1183)))},
                        $signed(wire1146)};
  assign wire1265 = $signed(reg1175);
  assign wire1266 = reg1173;
  always
    @(posedge clk) begin
      for (forvar1267 = (1'h0); (forvar1267 < (3'h4)); forvar1267 = (forvar1267 + (1'h1)))
        begin
          for (forvar1268 = (1'h0); (forvar1268 < (2'h3)); forvar1268 = (forvar1268 + (1'h1)))
            begin
              reg1269 <= ($signed({(|(reg1237 ? reg1164 : reg1237)),
                  $unsigned((reg1195 ?
                      wire1207 : reg1217))}) ^ (~^$signed($unsigned(reg1216))));
              reg1270 = ((+reg1160) & $unsigned(reg1237));
              reg1271 = (-{reg1270[(4'ha):(3'h5)]});
              reg1272 = (~|((reg1249[(4'h8):(3'h6)] ?
                      (8'hb9) : $unsigned(reg1183)) ?
                  (((reg1225 ? reg1198 : reg1216) ?
                      $unsigned((8'hab)) : $unsigned(reg1259)) * (+reg1153[(2'h2):(1'h0)])) : (&reg1220[(1'h0):(1'h0)])));
              reg1273 = reg1256[(1'h1):(1'h1)];
            end
          if ($signed($unsigned(wire1144)))
            begin
              reg1274 <= (reg1209 ^~ reg1222);
              reg1275 <= $unsigned($unsigned(reg1234[(4'hc):(1'h0)]));
              reg1276 = {(reg1271 ^ reg1203[(3'h5):(3'h4)])};
              reg1277 = (reg1200 ?
                  ((reg1248 ?
                      ({reg1194} ~^ $unsigned(reg1211)) : reg1249[(3'h4):(1'h0)]) == wire1207[(5'h16):(3'h7)]) : reg1234);
            end
          else
            begin
              reg1276 = $signed($unsigned($unsigned((wire1144[(4'h9):(1'h0)] && (~^reg1248)))));
              reg1277 = reg1237;
              reg1278 <= (~reg1184[(3'h6):(1'h1)]);
              reg1279 = $unsigned(($signed(($unsigned(reg1272) < (wire1264 ?
                  reg1168 : reg1160))) == $signed(reg1250[(5'h11):(5'h10)])));
              reg1280 <= ((reg1164[(1'h1):(1'h1)] * (((+reg1278) ?
                  (reg1234 << reg1175) : reg1253) | ($unsigned(reg1234) ?
                  $signed(reg1256) : $unsigned(reg1256)))) || (7'h42));
            end
          reg1281 <= wire1171[(3'h7):(2'h2)];
          reg1282 = wire1147[(4'h8):(2'h2)];
          if (wire1143[(3'h7):(3'h5)])
            begin
              reg1283 = (8'h9f);
            end
          else
            begin
              reg1283 = (|(~(~reg1273)));
              reg1284 <= $unsigned((+forvar1268));
            end
        end
      reg1285 <= reg1160;
      reg1286 = (reg1272[(4'ha):(1'h0)] <<< forvar1267);
      reg1287 = $unsigned($unsigned(reg1228));
    end
  always
    @(posedge clk) begin
      for (forvar1288 = (1'h0); (forvar1288 < (1'h1)); forvar1288 = (forvar1288 + (1'h1)))
        begin
          reg1289 = reg1205[(4'h9):(4'h9)];
        end
      reg1290 = $unsigned(reg1250);
      reg1291 <= $unsigned($unsigned($unsigned(((reg1158 ?
          wire1172 : reg1257) >> (reg1284 ? (8'h9e) : reg1211)))));
      for (forvar1292 = (1'h0); (forvar1292 < (2'h2)); forvar1292 = (forvar1292 + (1'h1)))
        begin
          if (($signed(reg1173[(5'h17):(2'h2)]) * {reg1228,
              (^(((8'ha5) | (8'hb7)) + reg1280))}))
            begin
              reg1293 <= ({$unsigned(((reg1278 ?
                          reg1184 : (8'ha9)) ^~ wire1148))} ?
                  {wire1144,
                      (|$signed(forvar1288[(3'h4):(2'h3)]))} : $unsigned((+(&((7'h40) ?
                      wire1207 : reg1194)))));
            end
          else
            begin
              reg1294 = reg1191[(3'h4):(2'h2)];
              reg1295 <= (reg1253[(2'h3):(2'h2)] ?
                  reg1218 : (~reg1249[(2'h2):(1'h1)]));
              reg1296 = ($unsigned((reg1151[(3'h6):(1'h0)] ?
                  reg1199 : reg1293)) >> wire1144);
            end
        end
      reg1297 <= ((reg1237 ?
          reg1184 : $unsigned(wire1146)) >>> {$signed(((reg1190 ?
                  reg1211 : (8'hb7)) ?
              reg1183[(3'h4):(2'h2)] : $signed(reg1293)))});
    end
  always
    @(posedge clk) begin
      for (forvar1298 = (1'h0); (forvar1298 < (1'h1)); forvar1298 = (forvar1298 + (1'h1)))
        begin
          reg1299 <= (reg1285 ?
              ((reg1173 ^ $unsigned({(8'ha9)})) ?
                  $unsigned((^$signed((8'haa)))) : (|((8'h9e) ?
                      (&wire1215) : reg1284[(4'hc):(3'h7)]))) : (^(~^reg1185)));
          reg1300 <= reg1256;
          reg1301 <= ((reg1195 >>> $unsigned(reg1293[(4'h8):(4'h8)])) ?
              $signed({reg1297}) : wire1171);
        end
      reg1302 = wire1143;
      for (forvar1303 = (1'h0); (forvar1303 < (2'h3)); forvar1303 = (forvar1303 + (1'h1)))
        begin
          if ((^~(7'h41)))
            begin
              reg1304 <= reg1173;
            end
          else
            begin
              reg1304 <= $unsigned((~^($signed(reg1300) ?
                  (^{reg1284, reg1256}) : ({(8'hab), reg1205} ?
                      (reg1302 ~^ reg1200) : (reg1300 ? reg1228 : reg1164)))));
              reg1305 <= ({{$unsigned((-wire1206)),
                          $signed({wire1144, (8'hae)})},
                      reg1191} ?
                  reg1208[(3'h4):(3'h4)] : ((+{reg1301}) ?
                      $signed(wire1147) : (|$signed((reg1195 << wire1266)))));
              reg1306 = $signed($unsigned($unsigned((8'haa))));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar1307 = (1'h0); (forvar1307 < (2'h3)); forvar1307 = (forvar1307 + (1'h1)))
        begin
          for (forvar1308 = (1'h0); (forvar1308 < (2'h3)); forvar1308 = (forvar1308 + (1'h1)))
            begin
              reg1309 <= reg1253;
              reg1310 = reg1175[(4'hd):(3'h7)];
              reg1311 = reg1297;
            end
          reg1312 = (($signed((^{(8'ha8), reg1299})) == $unsigned({(reg1185 ?
                      reg1256 : reg1164),
                  (reg1250 ? reg1284 : reg1183)})) ?
              ((~&{reg1281[(4'h9):(3'h6)]}) ?
                  reg1259[(4'h8):(1'h0)] : reg1281) : $signed(wire1143));
          reg1313 = (($unsigned(reg1223[(3'h5):(3'h5)]) ?
              $unsigned((+{(8'ha1), reg1185})) : $signed((((8'ha0) ?
                      reg1181 : reg1190) ?
                  (+reg1200) : $signed(wire1146)))) + wire1264[(4'hc):(3'h7)]);
          reg1314 <= $signed($signed($signed($unsigned(reg1151))));
          reg1315 = $unsigned((-{reg1257[(2'h3):(2'h2)], wire1264}));
        end
      reg1316 = $unsigned(wire1146);
      for (forvar1317 = (1'h0); (forvar1317 < (3'h4)); forvar1317 = (forvar1317 + (1'h1)))
        begin
          for (forvar1318 = (1'h0); (forvar1318 < (2'h2)); forvar1318 = (forvar1318 + (1'h1)))
            begin
              reg1319 = reg1300;
              reg1320 = reg1205[(2'h2):(1'h1)];
            end
          reg1321 <= {(wire1265 && ((&{(8'hb2)}) ?
                  (|(reg1269 && (7'h46))) : {reg1164}))};
          reg1322 = $unsigned((^~($signed((forvar1308 ^~ wire1207)) >= reg1153[(2'h3):(1'h0)])));
          for (forvar1323 = (1'h0); (forvar1323 < (1'h0)); forvar1323 = (forvar1323 + (1'h1)))
            begin
              reg1324 = ((({(reg1177 & (8'had))} ?
                  (8'hbe) : $unsigned($signed(reg1275))) & $signed($signed((~&reg1291)))) || reg1184[(3'h5):(3'h5)]);
              reg1325 <= reg1278[(4'hb):(4'ha)];
            end
        end
      for (forvar1326 = (1'h0); (forvar1326 < (2'h3)); forvar1326 = (forvar1326 + (1'h1)))
        begin
          reg1327 = (8'hba);
          reg1328 = {{reg1236[(1'h1):(1'h1)],
                  ($unsigned(((8'hbb) < wire1171)) ^ (reg1299[(4'hf):(3'h7)] ?
                      (+reg1181) : reg1291[(1'h0):(1'h0)]))},
              ({$unsigned((reg1300 <<< reg1259))} != (&((^reg1281) >>> reg1209[(1'h0):(1'h0)])))};
          for (forvar1329 = (1'h0); (forvar1329 < (1'h1)); forvar1329 = (forvar1329 + (1'h1)))
            begin
              reg1330 = (reg1229[(1'h1):(1'h0)] < {reg1259,
                  $unsigned((!$unsigned(reg1236)))});
              reg1331 <= (reg1179 ^~ reg1228);
              reg1332 <= ($signed(((reg1257 & {(8'hb3)}) ?
                      wire1143 : reg1228[(3'h5):(1'h0)])) ?
                  (7'h49) : {$unsigned({(reg1194 * reg1228)})});
              reg1333 <= (reg1281[(4'h8):(3'h4)] ?
                  reg1257[(3'h5):(1'h1)] : {$unsigned(reg1332[(2'h3):(2'h2)]),
                      {(((8'h9e) && wire1264) >> reg1236[(2'h3):(1'h1)]),
                          (~|{(8'had)})}});
              reg1334 = {reg1301, $signed(reg1209)};
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module937
#(parameter param1136 = (|{((((8'hb5) ? (8'hb2) : (8'hb5)) ? (!(8'ha2)) : (8'ha8)) ? ({(8'hb7)} ? ((7'h49) - (7'h4a)) : {(8'haa)}) : (8'hae)), {(((8'had) | (8'hb8)) || (~|(8'hae))), ({(8'h9d)} >>> ((8'hb6) > (8'haa)))}}), 
parameter param1137 = (~&param1136))
(y, clk, wire941, wire940, wire939, wire938);
  output wire [(32'ha0a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire941;
  input wire signed [(5'h14):(1'h0)] wire940;
  input wire [(4'h8):(1'h0)] wire939;
  input wire signed [(5'h17):(1'h0)] wire938;
  wire signed [(5'h13):(1'h0)] wire1131;
  wire [(4'ha):(1'h0)] wire1130;
  wire [(4'hf):(1'h0)] wire1129;
  wire [(5'h17):(1'h0)] wire1108;
  wire [(2'h2):(1'h0)] wire1060;
  wire signed [(5'h17):(1'h0)] wire1058;
  wire signed [(4'ha):(1'h0)] wire1057;
  wire [(3'h4):(1'h0)] wire1056;
  wire signed [(4'h8):(1'h0)] wire1055;
  wire signed [(5'h10):(1'h0)] wire1021;
  wire signed [(4'h8):(1'h0)] wire942;
  reg signed [(4'ha):(1'h0)] reg1134 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1132 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1126 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1122 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1121 = (1'h0);
  reg [(2'h3):(1'h0)] reg1120 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1117 = (1'h0);
  reg [(5'h15):(1'h0)] reg1112 = (1'h0);
  reg [(5'h13):(1'h0)] reg1110 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1107 = (1'h0);
  reg [(4'he):(1'h0)] reg1106 = (1'h0);
  reg [(5'h12):(1'h0)] reg1104 = (1'h0);
  reg [(2'h2):(1'h0)] reg1102 = (1'h0);
  reg [(5'h17):(1'h0)] reg1099 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1096 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1095 = (1'h0);
  reg [(5'h11):(1'h0)] reg1092 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1088 = (1'h0);
  reg [(5'h14):(1'h0)] reg1087 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1084 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1081 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1079 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1078 = (1'h0);
  reg [(4'hb):(1'h0)] reg1077 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1076 = (1'h0);
  reg [(4'hf):(1'h0)] reg1074 = (1'h0);
  reg [(5'h11):(1'h0)] reg1073 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1071 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1070 = (1'h0);
  reg [(3'h5):(1'h0)] reg1069 = (1'h0);
  reg [(4'hc):(1'h0)] reg1067 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1065 = (1'h0);
  reg [(4'ha):(1'h0)] reg1064 = (1'h0);
  reg [(5'h18):(1'h0)] reg1063 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1061 = (1'h0);
  reg [(4'hb):(1'h0)] reg1059 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1053 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1051 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1049 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1046 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1040 = (1'h0);
  reg [(4'h8):(1'h0)] reg1038 = (1'h0);
  reg [(4'ha):(1'h0)] reg1037 = (1'h0);
  reg [(3'h6):(1'h0)] reg1034 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1030 = (1'h0);
  reg [(5'h13):(1'h0)] reg1029 = (1'h0);
  reg [(3'h7):(1'h0)] reg1026 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1023 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1020 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1017 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1003 = (1'h0);
  reg [(5'h15):(1'h0)] reg1015 = (1'h0);
  reg [(3'h7):(1'h0)] reg1013 = (1'h0);
  reg [(5'h18):(1'h0)] reg1012 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1011 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1010 = (1'h0);
  reg [(4'hb):(1'h0)] reg1008 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1004 = (1'h0);
  reg [(4'hc):(1'h0)] reg1000 = (1'h0);
  reg [(4'hd):(1'h0)] reg998 = (1'h0);
  reg signed [(4'he):(1'h0)] reg996 = (1'h0);
  reg [(5'h18):(1'h0)] reg990 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg987 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg982 = (1'h0);
  reg [(3'h6):(1'h0)] reg980 = (1'h0);
  reg [(3'h5):(1'h0)] reg977 = (1'h0);
  reg [(2'h3):(1'h0)] reg974 = (1'h0);
  reg [(5'h10):(1'h0)] reg969 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg966 = (1'h0);
  reg [(5'h11):(1'h0)] reg964 = (1'h0);
  reg [(4'hf):(1'h0)] reg961 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg959 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg956 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg955 = (1'h0);
  reg [(4'hf):(1'h0)] reg954 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg949 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg947 = (1'h0);
  reg [(4'hb):(1'h0)] reg946 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg945 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1135 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1133 = (1'h0);
  reg [(5'h11):(1'h0)] reg1128 = (1'h0);
  reg [(5'h16):(1'h0)] reg1127 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1125 = (1'h0);
  reg [(5'h15):(1'h0)] reg1124 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1123 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1119 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1118 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1116 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1115 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1114 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1113 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1111 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1109 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1105 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1103 = (1'h0);
  reg [(3'h4):(1'h0)] forvar1101 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1100 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar1091 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1098 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1097 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1094 = (1'h0);
  reg [(3'h4):(1'h0)] reg1093 = (1'h0);
  reg [(4'hf):(1'h0)] reg1091 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1090 = (1'h0);
  reg [(4'h8):(1'h0)] reg1089 = (1'h0);
  reg [(2'h2):(1'h0)] reg1086 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1085 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1075 = (1'h0);
  reg [(4'ha):(1'h0)] reg1083 = (1'h0);
  reg [(4'hb):(1'h0)] reg1082 = (1'h0);
  reg [(5'h10):(1'h0)] reg1080 = (1'h0);
  reg [(4'h8):(1'h0)] reg1075 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1072 = (1'h0);
  reg [(5'h14):(1'h0)] reg1068 = (1'h0);
  reg [(5'h14):(1'h0)] reg1066 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1062 = (1'h0);
  reg [(4'hd):(1'h0)] reg1054 = (1'h0);
  reg [(5'h12):(1'h0)] reg1052 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1050 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1048 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1047 = (1'h0);
  reg [(3'h4):(1'h0)] reg1045 = (1'h0);
  reg [(3'h5):(1'h0)] reg1044 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1043 = (1'h0);
  reg [(4'he):(1'h0)] reg1042 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1041 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1039 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1036 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1035 = (1'h0);
  reg [(4'h8):(1'h0)] reg1033 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1032 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1031 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar1025 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1024 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1022 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1028 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1027 = (1'h0);
  reg [(5'h14):(1'h0)] reg1025 = (1'h0);
  reg [(4'h9):(1'h0)] forvar1024 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1022 = (1'h0);
  reg [(5'h11):(1'h0)] reg1019 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1018 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1007 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1016 = (1'h0);
  reg [(5'h11):(1'h0)] reg1014 = (1'h0);
  reg [(4'he):(1'h0)] reg1009 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1007 = (1'h0);
  reg [(5'h12):(1'h0)] reg1006 = (1'h0);
  reg [(5'h18):(1'h0)] reg1005 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1003 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1002 = (1'h0);
  reg [(2'h2):(1'h0)] reg1001 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg999 = (1'h0);
  reg [(5'h14):(1'h0)] forvar997 = (1'h0);
  reg [(4'hc):(1'h0)] reg997 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg995 = (1'h0);
  reg [(3'h5):(1'h0)] reg994 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg993 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg992 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar991 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar977 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg989 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg988 = (1'h0);
  reg [(5'h18):(1'h0)] reg986 = (1'h0);
  reg [(5'h11):(1'h0)] reg985 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg984 = (1'h0);
  reg [(4'hf):(1'h0)] reg983 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg981 = (1'h0);
  reg [(5'h13):(1'h0)] reg979 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg978 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg976 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar975 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg973 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg972 = (1'h0);
  reg [(4'he):(1'h0)] reg971 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg970 = (1'h0);
  reg [(5'h10):(1'h0)] forvar968 = (1'h0);
  reg [(2'h2):(1'h0)] reg967 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar965 = (1'h0);
  reg [(4'h8):(1'h0)] reg963 = (1'h0);
  reg [(5'h18):(1'h0)] reg962 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar960 = (1'h0);
  reg [(3'h5):(1'h0)] reg958 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg957 = (1'h0);
  reg [(4'h8):(1'h0)] forvar953 = (1'h0);
  reg [(4'hb):(1'h0)] reg952 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg951 = (1'h0);
  reg [(4'he):(1'h0)] reg950 = (1'h0);
  reg [(4'ha):(1'h0)] reg948 = (1'h0);
  reg [(2'h2):(1'h0)] reg944 = (1'h0);
  reg [(3'h4):(1'h0)] reg943 = (1'h0);
  assign y = {wire1131,
                 wire1130,
                 wire1129,
                 wire1108,
                 wire1060,
                 wire1058,
                 wire1057,
                 wire1056,
                 wire1055,
                 wire1021,
                 wire942,
                 reg1134,
                 reg1132,
                 reg1126,
                 reg1122,
                 reg1121,
                 reg1120,
                 reg1117,
                 reg1112,
                 reg1110,
                 reg1107,
                 reg1106,
                 reg1104,
                 reg1102,
                 reg1099,
                 reg1096,
                 reg1095,
                 reg1092,
                 reg1088,
                 reg1087,
                 reg1084,
                 reg1081,
                 reg1079,
                 reg1078,
                 reg1077,
                 reg1076,
                 reg1074,
                 reg1073,
                 reg1071,
                 reg1070,
                 reg1069,
                 reg1067,
                 reg1065,
                 reg1064,
                 reg1063,
                 reg1061,
                 reg1059,
                 reg1053,
                 reg1051,
                 reg1049,
                 reg1046,
                 reg1040,
                 reg1038,
                 reg1037,
                 reg1034,
                 reg1030,
                 reg1029,
                 reg1026,
                 reg1023,
                 reg1020,
                 reg1017,
                 reg1003,
                 reg1015,
                 reg1013,
                 reg1012,
                 reg1011,
                 reg1010,
                 reg1008,
                 reg1004,
                 reg1000,
                 reg998,
                 reg996,
                 reg990,
                 reg987,
                 reg982,
                 reg980,
                 reg977,
                 reg974,
                 reg969,
                 reg966,
                 reg964,
                 reg961,
                 reg959,
                 reg956,
                 reg955,
                 reg954,
                 reg949,
                 reg947,
                 reg946,
                 reg945,
                 reg1135,
                 forvar1133,
                 reg1128,
                 reg1127,
                 forvar1125,
                 reg1124,
                 forvar1123,
                 forvar1119,
                 reg1118,
                 reg1116,
                 reg1115,
                 forvar1114,
                 reg1113,
                 forvar1111,
                 forvar1109,
                 reg1105,
                 reg1103,
                 forvar1101,
                 reg1100,
                 forvar1091,
                 reg1098,
                 reg1097,
                 reg1094,
                 reg1093,
                 reg1091,
                 reg1090,
                 reg1089,
                 reg1086,
                 forvar1085,
                 forvar1075,
                 reg1083,
                 reg1082,
                 reg1080,
                 reg1075,
                 reg1072,
                 reg1068,
                 reg1066,
                 reg1062,
                 reg1054,
                 reg1052,
                 forvar1050,
                 reg1048,
                 reg1047,
                 reg1045,
                 reg1044,
                 forvar1043,
                 reg1042,
                 forvar1041,
                 reg1039,
                 reg1036,
                 reg1035,
                 reg1033,
                 forvar1032,
                 reg1031,
                 forvar1025,
                 reg1024,
                 reg1022,
                 reg1028,
                 reg1027,
                 reg1025,
                 forvar1024,
                 forvar1022,
                 reg1019,
                 reg1018,
                 reg1007,
                 reg1016,
                 reg1014,
                 reg1009,
                 forvar1007,
                 reg1006,
                 reg1005,
                 forvar1003,
                 reg1002,
                 reg1001,
                 reg999,
                 forvar997,
                 reg997,
                 reg995,
                 reg994,
                 reg993,
                 reg992,
                 forvar991,
                 forvar977,
                 reg989,
                 reg988,
                 reg986,
                 reg985,
                 reg984,
                 reg983,
                 reg981,
                 reg979,
                 reg978,
                 reg976,
                 forvar975,
                 reg973,
                 reg972,
                 reg971,
                 reg970,
                 forvar968,
                 reg967,
                 forvar965,
                 reg963,
                 reg962,
                 forvar960,
                 reg958,
                 reg957,
                 forvar953,
                 reg952,
                 reg951,
                 reg950,
                 reg948,
                 reg944,
                 reg943,
                 (1'h0)};
  assign wire942 = (8'ha8);
  always
    @(posedge clk) begin
      if ((~|(wire942[(4'h8):(3'h6)] ^~ $unsigned((wire941 ?
          wire939[(4'h8):(3'h4)] : (wire942 ? wire942 : wire941))))))
        begin
          reg943 = wire939[(3'h4):(1'h0)];
          reg944 = wire942[(3'h6):(3'h5)];
          reg945 <= $signed(wire938);
        end
      else
        begin
          if ($unsigned(($signed((+(wire940 < wire938))) ?
              {((^wire938) <= reg944),
                  ((reg943 ? reg945 : (8'hb1)) ?
                      (reg944 ?
                          reg943 : (8'hbf)) : $signed(wire942))} : wire941)))
            begin
              reg945 <= (wire938 * ($unsigned(((7'h4a) <= (~|wire938))) ?
                  (~&wire940[(2'h2):(2'h2)]) : {wire938[(4'hf):(4'he)]}));
              reg946 <= wire940[(1'h0):(1'h0)];
              reg947 <= $unsigned((!wire940[(3'h6):(3'h4)]));
              reg948 = reg947[(4'h9):(3'h4)];
              reg949 <= wire941[(4'hd):(3'h5)];
            end
          else
            begin
              reg945 <= (|reg945[(2'h2):(1'h0)]);
              reg948 = reg948;
              reg950 = wire942[(3'h6):(3'h4)];
              reg951 = $unsigned((~|wire939));
              reg952 = reg943[(2'h3):(2'h2)];
            end
          for (forvar953 = (1'h0); (forvar953 < (3'h4)); forvar953 = (forvar953 + (1'h1)))
            begin
              reg954 <= reg950;
              reg955 <= ((($signed($unsigned(wire942)) ?
                  ($signed(wire938) ?
                      $signed(reg951) : (~|wire938)) : (wire942[(1'h1):(1'h0)] < $unsigned(wire941))) + ((8'h9d) ?
                  $signed({wire938}) : $unsigned(wire940))) >>> $signed((8'hba)));
              reg956 <= (|reg946[(2'h2):(1'h1)]);
              reg957 = $signed($signed((((reg952 && (8'ha3)) ?
                      $signed(wire939) : (reg945 ? reg946 : reg954)) ?
                  $signed(reg956) : $unsigned($unsigned(reg949)))));
            end
          reg958 = wire940[(3'h5):(3'h5)];
          reg959 <= {$unsigned($signed(reg955)), reg945};
          for (forvar960 = (1'h0); (forvar960 < (2'h2)); forvar960 = (forvar960 + (1'h1)))
            begin
              reg961 <= (|(^$unsigned(($signed((8'haa)) ?
                  $unsigned(reg958) : (reg945 ? reg943 : reg950)))));
              reg962 = (^~(reg946[(3'h5):(3'h4)] ?
                  $unsigned($unsigned((reg957 >>> reg959))) : $signed((8'haf))));
              reg963 = wire938;
              reg964 <= reg963;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar965 = (1'h0); (forvar965 < (1'h0)); forvar965 = (forvar965 + (1'h1)))
        begin
          reg966 <= (wire940[(3'h6):(3'h4)] ?
              ($unsigned((wire941[(4'hd):(3'h4)] ?
                      $unsigned(wire941) : $signed(reg949))) ?
                  ($signed($signed(reg947)) ?
                      {$unsigned(reg949)} : ($signed(reg949) * (reg964 ?
                          wire938 : (7'h43)))) : (-{(reg945 <= reg946)})) : wire940);
          reg967 = reg966[(1'h1):(1'h1)];
          for (forvar968 = (1'h0); (forvar968 < (1'h1)); forvar968 = (forvar968 + (1'h1)))
            begin
              reg969 <= (reg946 ?
                  ($unsigned(({reg967} ?
                      (reg964 >= reg954) : (reg964 ?
                          reg946 : wire942))) && $unsigned({reg964[(2'h2):(1'h0)],
                      {(8'h9c), (8'ha1)}})) : (-{wire938, (!(^wire941))}));
              reg970 = {wire939[(3'h6):(3'h4)], (^reg967[(2'h2):(1'h1)])};
              reg971 = $unsigned(((reg956[(4'hb):(3'h7)] ?
                      (~reg961[(2'h3):(2'h3)]) : reg969) ?
                  $signed((&wire942)) : (((|reg961) ?
                          (forvar968 ? (8'h9c) : reg945) : reg964) ?
                      reg946 : $unsigned((~reg949)))));
              reg972 = wire940[(3'h7):(3'h7)];
              reg973 = (^~$unsigned({$signed(wire939), wire941}));
            end
          reg974 <= wire941[(4'he):(1'h1)];
          for (forvar975 = (1'h0); (forvar975 < (3'h4)); forvar975 = (forvar975 + (1'h1)))
            begin
              reg976 = (8'hb6);
            end
        end
      if (((((^~(reg972 ? (7'h49) : wire938)) >>> $unsigned((reg974 ?
              reg949 : reg976))) >> ({$unsigned(reg974)} ?
              (&(8'ha4)) : ((reg956 ?
                  (8'hb4) : reg966) << $unsigned(reg970)))) ?
          reg972 : (({reg947, $signed(reg973)} ?
                  ($unsigned(forvar965) ?
                      ((8'hb4) ?
                          reg954 : reg947) : (!wire941)) : $unsigned($unsigned(reg949))) ?
              $unsigned(reg945[(3'h5):(1'h1)]) : $unsigned(wire942))))
        begin
          if ($unsigned((^$unsigned((reg970[(5'h13):(4'hd)] ?
              wire938 : $signed(wire939))))))
            begin
              reg977 <= ($unsigned((reg967 ?
                      (^~(8'hbf)) : (reg945[(2'h2):(1'h0)] ?
                          reg955[(3'h5):(2'h3)] : reg966))) ?
                  reg959[(3'h5):(3'h4)] : {$signed(reg945)});
              reg978 = reg973;
              reg979 = $signed(({((reg978 >= reg966) && reg977[(1'h0):(1'h0)])} ?
                  $signed(reg959[(1'h1):(1'h1)]) : reg969));
              reg980 <= ($unsigned((($signed(reg947) - (wire942 ?
                      reg945 : forvar975)) ?
                  {$unsigned(reg977)} : {forvar975[(5'h10):(4'hf)],
                      $signed(reg971)})) * (forvar975[(4'h9):(3'h5)] ?
                  ($signed((wire939 ? reg970 : (8'ha5))) || ((reg970 ?
                      wire940 : forvar975) ~^ (reg961 ?
                      reg972 : reg967))) : ($unsigned($signed((7'h40))) >= ((wire938 ?
                          wire940 : reg964) ?
                      $unsigned((8'hb2)) : (reg966 > reg977)))));
              reg981 = reg974;
            end
          else
            begin
              reg978 = reg978[(2'h2):(1'h1)];
              reg979 = (&forvar968);
              reg980 <= (^~$unsigned($signed($signed((~&(7'h40))))));
              reg982 <= reg961[(4'ha):(3'h5)];
              reg983 = reg977;
            end
          reg984 = $unsigned(reg955);
          reg985 = (~|$unsigned(reg969[(3'h4):(2'h2)]));
          reg986 = $signed($unsigned($unsigned(reg976[(3'h7):(3'h5)])));
          if ($signed(((~|(^~reg979[(4'hf):(4'h8)])) ~^ $signed(reg947))))
            begin
              reg987 <= $signed($unsigned((($unsigned(reg956) ?
                      ((8'hb3) == (8'ha6)) : wire941[(4'h9):(3'h4)]) ?
                  $unsigned($unsigned(reg973)) : ($signed((8'hb7)) ?
                      $signed(reg984) : reg979))));
              reg988 = $signed(reg976);
              reg989 = (reg954[(4'hd):(4'h8)] ?
                  (reg983[(4'he):(3'h5)] ?
                      $signed(reg969[(5'h10):(3'h5)]) : reg983[(4'hb):(4'hb)]) : (reg955 ?
                      $unsigned(reg978[(1'h1):(1'h0)]) : (forvar968[(4'hb):(4'hb)] & (reg983[(2'h2):(1'h1)] ?
                          $signed(reg961) : (~^(7'h44))))));
            end
          else
            begin
              reg987 <= ({($unsigned({reg966,
                      reg986}) >>> reg974[(1'h0):(1'h0)]),
                  {({reg959, reg985} ?
                          (reg949 ? (7'h46) : reg947) : (~^reg988)),
                      reg966}} + (~&({$signed(reg976)} ~^ (!$unsigned(wire938)))));
              reg988 = (~&(reg961[(3'h5):(3'h5)] ?
                  $signed(reg988[(4'hb):(3'h5)]) : $signed(({reg954} < {reg973}))));
              reg990 <= $signed(reg970[(4'h8):(4'h8)]);
            end
        end
      else
        begin
          for (forvar977 = (1'h0); (forvar977 < (2'h2)); forvar977 = (forvar977 + (1'h1)))
            begin
              reg980 <= (&({({reg980, reg973} && $unsigned((8'ha2))),
                  ((8'h9f) + $signed((8'h9f)))} >= {(((8'hbd) << reg969) ?
                      (reg980 >>> reg982) : reg954),
                  ($signed(reg986) || (reg987 * reg949))}));
              reg982 <= reg972[(4'hb):(1'h1)];
            end
          if (reg983)
            begin
              reg983 = wire942[(3'h7):(3'h7)];
              reg987 <= reg989;
              reg988 = (8'hb0);
              reg989 = $signed($signed($signed(reg947[(5'h10):(2'h3)])));
            end
          else
            begin
              reg983 = ((~((((8'hbe) | reg988) ?
                      (&reg988) : $unsigned(reg985)) ?
                  (reg970 ?
                      $signed(reg989) : $signed(reg954)) : $signed(((8'ha0) ?
                      (7'h41) : forvar975)))) + ($unsigned($unsigned((reg985 ?
                      (7'h4a) : reg977))) ?
                  wire942 : reg989));
              reg984 = $signed({(+($signed(reg976) ?
                      $signed(reg949) : reg972))});
              reg987 <= (((&(^~$signed(reg961))) == ((reg959[(4'h9):(4'h8)] ?
                      (~&reg959) : (reg981 ~^ forvar965)) ?
                  {{reg964}} : $signed($unsigned(reg959)))) + wire941);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar991 = (1'h0); (forvar991 < (1'h0)); forvar991 = (forvar991 + (1'h1)))
        begin
          reg992 = (|($signed($signed($unsigned(reg947))) ?
              ($signed($unsigned(wire939)) < $signed((wire942 <<< reg961))) : ($signed(reg980[(2'h3):(2'h3)]) != ((reg961 ^ forvar991) ?
                  $unsigned(wire941) : {reg956}))));
          reg993 = $signed((($signed((reg955 ? wire939 : reg974)) ?
                  ((~^(7'h46)) >= (-reg954)) : reg966) ?
              $signed((reg992[(4'hd):(4'h8)] ?
                  reg990 : (reg977 || (8'hae)))) : wire939));
          reg994 = $signed(reg961);
          reg995 = {(reg964[(4'h9):(3'h4)] ^~ {reg990[(4'h9):(3'h4)]}),
              $signed((!($signed((8'hb0)) ?
                  $signed(reg966) : (reg947 ~^ wire940))))};
          reg996 <= (($unsigned(((reg977 ? reg992 : (8'ha1)) ?
                  (^(8'ha6)) : (+reg992))) ~^ reg946) ?
              (reg954 ?
                  ($unsigned(reg945[(1'h0):(1'h0)]) ?
                      reg945[(2'h3):(1'h1)] : (!reg993)) : reg964) : (~^forvar991[(4'hc):(3'h5)]));
        end
      if ($unsigned(reg966))
        begin
          reg997 = ((reg992[(1'h1):(1'h1)] >> $signed(reg955[(3'h6):(2'h3)])) ?
              reg987 : ((reg995[(5'h10):(4'hb)] >>> reg982[(3'h6):(3'h5)]) >= (8'ha2)));
          reg998 <= (&(reg964[(4'hd):(3'h5)] && $unsigned($unsigned((reg956 ?
              (7'h43) : reg997)))));
        end
      else
        begin
          for (forvar997 = (1'h0); (forvar997 < (1'h0)); forvar997 = (forvar997 + (1'h1)))
            begin
              reg998 <= $unsigned(((reg996 ?
                  {reg996[(3'h6):(2'h3)]} : (-(reg992 ?
                      reg980 : reg987))) >> {$signed(((8'ha0) ?
                      reg946 : wire941)),
                  ($unsigned(reg974) ? (!reg969) : (~^reg990))}));
              reg999 = wire938;
              reg1000 <= (^$signed(reg955[(1'h1):(1'h1)]));
              reg1001 = reg959[(3'h6):(1'h1)];
            end
        end
      if ($unsigned((^~(~&(reg949 >>> (8'hbb))))))
        begin
          reg1002 = ((((^{reg974}) ?
              reg945 : (|(&reg945))) && (~^reg1001)) ^ $signed((~^{$unsigned((8'hab)),
              $signed((8'ha2))})));
          for (forvar1003 = (1'h0); (forvar1003 < (1'h0)); forvar1003 = (forvar1003 + (1'h1)))
            begin
              reg1004 <= (+$unsigned($unsigned((reg977[(3'h4):(3'h4)] ?
                  (-reg990) : $unsigned(reg947)))));
              reg1005 = $unsigned($signed(wire940));
              reg1006 = $unsigned($signed(reg995));
            end
          for (forvar1007 = (1'h0); (forvar1007 < (2'h3)); forvar1007 = (forvar1007 + (1'h1)))
            begin
              reg1008 <= $unsigned((|(!$unsigned($unsigned(reg947)))));
              reg1009 = $unsigned($unsigned($unsigned((!$signed(reg946)))));
              reg1010 <= (reg974 ?
                  (reg992[(5'h12):(1'h0)] ?
                      $signed({{reg961}}) : reg999[(1'h1):(1'h1)]) : ((((~^wire938) ?
                          (wire942 <= reg1004) : $signed(reg961)) ?
                      $unsigned(wire939) : $unsigned((reg1009 ?
                          reg947 : (8'hbe)))) >= reg949));
            end
          if ((~|reg945))
            begin
              reg1011 <= (!wire942);
              reg1012 <= ($unsigned(((7'h48) ? forvar997 : (~&(-(8'ha4))))) ?
                  ($signed((-(~reg947))) >>> $unsigned(($unsigned(reg946) ?
                      (forvar1007 ?
                          reg1001 : reg949) : reg1005[(4'hd):(3'h7)]))) : $unsigned($unsigned((+(reg954 ?
                      reg1002 : reg1011)))));
              reg1013 <= {$signed((~^((~&(7'h4a)) ?
                      (reg996 - reg982) : {reg999})))};
              reg1014 = ($unsigned(($signed($signed(reg997)) ?
                      $signed((reg1010 ?
                          reg966 : reg1010)) : {reg1011[(4'hd):(4'hb)],
                          (reg1002 >>> reg994)})) ?
                  reg1001[(1'h1):(1'h0)] : ((!wire941[(4'he):(4'he)]) ^~ ((^~$unsigned(reg1002)) >>> (~|$unsigned(wire942)))));
              reg1015 <= $unsigned($signed((($signed(reg993) == $signed(reg1011)) ?
                  (reg982 ?
                      $unsigned(reg947) : reg1006) : (reg1009[(4'hb):(4'hb)] ?
                      (reg993 ? reg947 : reg1004) : (reg993 >> reg966)))));
            end
          else
            begin
              reg1011 <= reg969;
            end
          reg1016 = $unsigned(((((reg974 ~^ forvar991) ?
              (reg966 ?
                  reg949 : reg1015) : $unsigned(forvar1003)) << $unsigned((|reg992))) ~^ (7'h44)));
        end
      else
        begin
          reg1002 = $unsigned($unsigned($signed(reg1014)));
          reg1003 <= ({$unsigned(($signed((7'h47)) ^~ wire940[(3'h6):(2'h2)])),
              reg977} ^~ $unsigned($unsigned(reg1002)));
          reg1005 = $unsigned($unsigned($unsigned((~|reg947[(1'h1):(1'h1)]))));
          reg1006 = reg995[(4'ha):(1'h1)];
          reg1007 = $unsigned($signed((~$unsigned((wire941 & reg1013)))));
        end
      reg1017 <= reg949[(4'h9):(1'h0)];
      if ($unsigned($signed($unsigned($unsigned((~^reg994))))))
        begin
          reg1018 = $signed($signed(reg1000));
          if ((&(8'hab)))
            begin
              reg1019 = $signed(($signed($signed($unsigned(reg969))) ?
                  (reg1002[(2'h3):(1'h0)] ?
                      (~|$unsigned(reg1012)) : $unsigned((forvar1007 + wire939))) : reg1014[(4'hf):(3'h5)]));
              reg1020 <= {(^reg998), reg1003[(1'h1):(1'h1)]};
            end
          else
            begin
              reg1020 <= ($unsigned((((+(8'hb9)) < {reg954}) ?
                  {(reg1000 ?
                          reg987 : forvar997)} : reg961)) <<< $unsigned(reg956[(5'h12):(2'h3)]));
            end
        end
      else
        begin
          reg1018 = ((&forvar1007[(1'h1):(1'h1)]) ?
              $signed(reg977) : $unsigned((~^reg1009)));
        end
    end
  assign wire1021 = (reg947[(5'h10):(4'hc)] ?
                        $unsigned($signed(((7'h42) < $signed((8'hbf))))) : $signed(((((8'ha0) ?
                            reg954 : reg954) ^ (~^reg977)) == (reg945 - reg982))));
  always
    @(posedge clk) begin
      if ((8'ha9))
        begin
          for (forvar1022 = (1'h0); (forvar1022 < (1'h0)); forvar1022 = (forvar1022 + (1'h1)))
            begin
              reg1023 <= (8'ha8);
            end
          for (forvar1024 = (1'h0); (forvar1024 < (2'h3)); forvar1024 = (forvar1024 + (1'h1)))
            begin
              reg1025 = $unsigned(reg1023);
              reg1026 <= $unsigned((reg1004 > (forvar1022[(3'h4):(1'h0)] ^~ reg974[(1'h1):(1'h1)])));
              reg1027 = reg1020;
              reg1028 = (wire938[(5'h15):(5'h11)] != ($unsigned(reg969) ?
                  ((~&reg1017) >>> ($signed(reg969) ?
                      $unsigned(reg1011) : reg1017[(3'h4):(2'h2)])) : ($unsigned(reg980) >> $signed((~&reg954)))));
            end
        end
      else
        begin
          reg1022 = (((7'h49) ?
                  (~|((reg990 ?
                      (8'ha8) : reg990) & reg1028[(4'h8):(4'h8)])) : $signed((reg969[(4'hf):(1'h1)] <<< (reg955 ?
                      reg961 : reg977)))) ?
              {(reg954 != {(!reg1017)})} : (&(-reg1010[(4'hc):(3'h4)])));
          reg1024 = (($unsigned((!reg1017[(3'h5):(3'h5)])) ?
              $signed((|(-(8'hbc)))) : reg1017[(2'h3):(2'h3)]) > reg977);
          for (forvar1025 = (1'h0); (forvar1025 < (1'h1)); forvar1025 = (forvar1025 + (1'h1)))
            begin
              reg1026 <= $signed($signed(($signed($unsigned(wire940)) ?
                  $unsigned($unsigned(reg947)) : (~$signed(reg1015)))));
              reg1029 <= $signed({$unsigned(wire938[(1'h1):(1'h1)])});
              reg1030 <= ($unsigned((reg949 ?
                      $unsigned($signed(reg945)) : ($signed(reg1010) & $unsigned(reg998)))) ?
                  (reg949 * $unsigned(forvar1022)) : $signed((~&reg961)));
            end
        end
      reg1031 = reg996[(3'h5):(1'h0)];
      for (forvar1032 = (1'h0); (forvar1032 < (1'h0)); forvar1032 = (forvar1032 + (1'h1)))
        begin
          reg1033 = (({((wire938 ^ (8'hbf)) ?
                      $unsigned(reg964) : ((8'hb6) << forvar1025))} & (^reg1012[(3'h5):(1'h1)])) ?
              (((reg955 <<< (reg1024 ?
                  reg1026 : wire938)) == ((reg955 == forvar1025) ?
                  $signed(reg1004) : (!forvar1032))) * $signed(reg987)) : reg949);
          reg1034 <= (~reg1031[(1'h0):(1'h0)]);
          reg1035 = ((^~$unsigned($signed((reg966 ? wire942 : reg1008)))) ?
              (8'hb7) : $unsigned($signed(wire938)));
          if (reg1031[(4'h8):(2'h2)])
            begin
              reg1036 = (~&(($signed($signed(wire940)) & {$signed(reg974),
                      $signed(reg977)}) ?
                  $unsigned(($signed((8'hb5)) && (forvar1025 < reg1029))) : $unsigned(reg1020[(1'h1):(1'h0)])));
              reg1037 <= ((~|$signed(reg974)) >> (!(&((wire941 ?
                      reg1022 : wire939) ?
                  $unsigned(reg982) : (reg1011 > reg1030)))));
              reg1038 <= {{{reg955[(1'h0):(1'h0)]},
                      $unsigned({(reg956 & reg1028)})},
                  (7'h44)};
            end
          else
            begin
              reg1037 <= reg990[(5'h16):(3'h4)];
              reg1038 <= reg982[(4'hd):(4'ha)];
              reg1039 = $unsigned($signed($signed($unsigned({(8'hb7),
                  reg959}))));
              reg1040 <= (!reg961[(4'he):(3'h6)]);
            end
          for (forvar1041 = (1'h0); (forvar1041 < (1'h0)); forvar1041 = (forvar1041 + (1'h1)))
            begin
              reg1042 = (((7'h42) || (&(8'hba))) ^~ $signed(($unsigned((reg1028 ^ reg1000)) != $unsigned($unsigned((8'hae))))));
            end
        end
      for (forvar1043 = (1'h0); (forvar1043 < (2'h2)); forvar1043 = (forvar1043 + (1'h1)))
        begin
          if ($signed(($unsigned($signed($signed(wire938))) << (7'h49))))
            begin
              reg1044 = wire940[(4'hb):(3'h6)];
              reg1045 = $signed({$unsigned(reg947[(5'h10):(4'ha)]),
                  $signed($unsigned((reg1036 >> reg947)))});
              reg1046 <= $signed($signed($signed(((+reg947) ~^ (reg1011 ?
                  (7'h43) : reg1012)))));
              reg1047 = {wire941,
                  ((+$unsigned((reg1013 ? reg1017 : reg959))) ?
                      (~reg961) : reg987[(3'h6):(3'h6)])};
            end
          else
            begin
              reg1046 <= reg969;
            end
          reg1048 = reg1013;
          reg1049 <= reg945[(3'h4):(3'h4)];
          for (forvar1050 = (1'h0); (forvar1050 < (2'h3)); forvar1050 = (forvar1050 + (1'h1)))
            begin
              reg1051 <= (~(-reg949));
              reg1052 = $unsigned($unsigned($unsigned((~&(wire939 ?
                  reg990 : reg974)))));
              reg1053 <= (^wire942);
              reg1054 = ({$unsigned(reg955)} > ($signed($unsigned({reg1031})) ^ {(^~{reg1036,
                      reg1017})}));
            end
        end
    end
  assign wire1055 = reg1037;
  assign wire1056 = (~&(^~reg1020));
  assign wire1057 = (&$signed((((wire939 ? reg1000 : reg956) ?
                        (~|reg998) : {reg980}) * $signed(reg1008))));
  assign wire1058 = wire942[(2'h3):(1'h0)];
  always
    @(posedge clk) begin
      reg1059 <= {reg987[(4'hf):(2'h3)]};
    end
  assign wire1060 = ((($unsigned((+(8'hbd))) || reg1038[(3'h7):(2'h3)]) >>> reg1030[(2'h2):(1'h0)]) ?
                        reg1034[(3'h4):(2'h3)] : ((($unsigned((7'h48)) ?
                                {reg1034} : wire1058[(3'h5):(2'h2)]) ?
                            (^$signed(reg998)) : (reg987[(4'hb):(3'h7)] ~^ (wire942 * reg1051))) ^ reg1037[(2'h2):(1'h0)]));
  always
    @(posedge clk) begin
      reg1061 <= (reg1010[(1'h0):(1'h0)] ^~ {(~((~^reg977) == (reg977 < (8'hb8))))});
      if ((~^reg1040))
        begin
          reg1062 = $signed(reg1061);
          if ((reg1037 >> {$unsigned($unsigned({reg977}))}))
            begin
              reg1063 <= (((~&{{(8'haf)},
                      reg982[(5'h13):(1'h0)]}) >>> ($signed(reg955) ?
                      (reg1034[(2'h3):(1'h1)] <<< (reg954 >> reg1037)) : $signed((wire939 * reg949)))) ?
                  (wire942 ?
                      $unsigned((&wire1056)) : reg996[(3'h5):(3'h5)]) : {((reg959 ?
                          wire939 : reg1049[(4'h8):(3'h5)]) >> $signed($unsigned((8'hbe))))});
              reg1064 <= (reg1046[(1'h0):(1'h0)] << (reg987[(5'h18):(4'he)] && ((wire1060[(2'h2):(2'h2)] & (reg1012 ?
                  reg996 : reg1013)) && ($signed(wire938) ?
                  (reg1020 ? reg1000 : wire940) : (8'hb2)))));
              reg1065 <= ($unsigned(($signed((reg998 ~^ reg1026)) ?
                  (reg1049 ? $unsigned(reg1063) : reg1011) : ((^wire1060) ?
                      ((7'h46) ?
                          (8'hb6) : reg990) : (reg1015 ^ reg1011)))) <= ((^~$unsigned(reg1061[(5'h13):(3'h4)])) >> reg969));
              reg1066 = (^$signed((((reg1062 ?
                  reg990 : reg946) <= (reg1062 || reg1037)) - $unsigned((reg1003 ?
                  reg980 : wire1021)))));
            end
          else
            begin
              reg1066 = {reg974,
                  ((&$signed((+reg1059))) ? (+{$signed(reg1008)}) : reg969)};
              reg1067 <= ((8'h9d) | $unsigned($signed((~|$unsigned(reg945)))));
              reg1068 = (reg1010[(4'hb):(2'h2)] >> (reg1034 ?
                  $signed($signed(reg1063[(4'hc):(3'h4)])) : {(|reg977[(3'h5):(1'h1)]),
                      reg955[(3'h4):(1'h0)]}));
            end
          if ($unsigned(reg1000))
            begin
              reg1069 <= $signed((^~$signed($signed($signed(wire939)))));
              reg1070 <= (((wire1021[(3'h4):(1'h0)] >>> (~(reg945 | reg1059))) >> (reg1030 << $unsigned({reg1065}))) + $unsigned(reg945));
              reg1071 <= {reg1064[(3'h5):(1'h0)]};
            end
          else
            begin
              reg1072 = $unsigned($signed((8'hbf)));
              reg1073 <= (reg998[(2'h2):(1'h0)] != reg954[(3'h7):(1'h1)]);
            end
        end
      else
        begin
          reg1062 = $signed(reg946[(4'hb):(3'h4)]);
        end
      reg1074 <= {$signed((($signed((8'h9e)) - (!reg964)) ?
              reg945 : ((!reg1051) || wire1057[(3'h6):(3'h5)])))};
    end
  always
    @(posedge clk) begin
      if ($unsigned($unsigned($unsigned((reg949 ~^ $unsigned(reg956))))))
        begin
          reg1075 = ($unsigned($unsigned(reg1053[(1'h1):(1'h1)])) >>> reg966);
          reg1076 <= {$signed(wire941[(3'h4):(2'h3)])};
          reg1077 <= wire938;
          reg1078 <= reg969;
          if (((|(~&((reg1004 < reg1049) ?
              ((7'h46) << (8'haa)) : $unsigned(reg1017)))) > (($signed((+(8'ha0))) <<< $signed(reg974[(1'h1):(1'h0)])) ?
              $unsigned(((reg1064 ? reg966 : reg1075) ?
                  reg1069[(2'h3):(2'h3)] : reg1008[(4'ha):(4'ha)])) : $unsigned($signed((reg1011 ?
                  reg1023 : reg964))))))
            begin
              reg1079 <= ((reg961 ?
                      (-(reg998 * (^reg1040))) : ($signed(reg1003[(5'h11):(3'h6)]) ?
                          wire939 : ($unsigned(reg1010) ^ $unsigned(reg1034)))) ?
                  (wire1021[(4'h8):(1'h1)] ?
                      $unsigned($signed(reg1069)) : ((^~wire1058[(5'h15):(5'h14)]) ?
                          (8'ha5) : (8'hbc))) : $signed(($unsigned((!(8'hb7))) ?
                      (wire938 <<< (reg1020 ?
                          (7'h42) : (7'h47))) : reg959[(1'h0):(1'h0)])));
              reg1080 = $unsigned(reg956);
              reg1081 <= $unsigned(reg946);
              reg1082 = ({reg1071[(3'h5):(1'h1)]} + (reg1012[(4'h9):(3'h7)] * (reg1049 ?
                  (|reg1079[(4'h8):(3'h7)]) : reg1078[(1'h1):(1'h0)])));
              reg1083 = $unsigned({{reg1029}});
            end
          else
            begin
              reg1080 = (~|$signed(wire1056[(2'h2):(1'h1)]));
              reg1081 <= (&$unsigned(reg1023[(2'h3):(2'h3)]));
            end
        end
      else
        begin
          for (forvar1075 = (1'h0); (forvar1075 < (3'h4)); forvar1075 = (forvar1075 + (1'h1)))
            begin
              reg1076 <= reg998[(4'ha):(4'ha)];
              reg1080 = $signed((wire1055[(3'h4):(1'h1)] ?
                  (~$unsigned((~|reg974))) : (^~$unsigned($unsigned((8'hb9))))));
              reg1081 <= (reg954 < (~(~|$unsigned(reg966))));
              reg1084 <= ((reg977 ?
                  $signed(forvar1075[(3'h7):(1'h1)]) : $unsigned((-$unsigned(reg961)))) != (!{{reg1046,
                      reg1076[(3'h6):(1'h1)]}}));
            end
          for (forvar1085 = (1'h0); (forvar1085 < (3'h4)); forvar1085 = (forvar1085 + (1'h1)))
            begin
              reg1086 = ($unsigned((~&reg947[(1'h1):(1'h0)])) ?
                  $signed(((&$signed(reg998)) ?
                      $signed((8'hab)) : $signed((-(8'hbf))))) : ($signed(($signed(reg969) ?
                          (wire942 && reg1017) : (~&reg1017))) ?
                      reg1008[(2'h3):(2'h3)] : (reg959 * $signed(reg1083[(4'h8):(4'h8)]))));
            end
          reg1087 <= {reg980[(2'h3):(2'h3)]};
          reg1088 <= reg1015;
        end
      reg1089 = {$signed($unsigned((~&$signed(reg1087))))};
      if (reg1010)
        begin
          reg1090 = $unsigned(reg1034[(3'h4):(2'h2)]);
          reg1091 = $unsigned((&reg1087));
          if ($unsigned({$unsigned(reg1087)}))
            begin
              reg1092 <= (&(~^$unsigned((^~(!(8'hb6))))));
              reg1093 = $unsigned((($signed(reg1070[(2'h2):(2'h2)]) ?
                      reg1082[(1'h1):(1'h1)] : wire1021) ?
                  reg1017 : (^reg1089[(3'h6):(1'h0)])));
              reg1094 = reg1023;
              reg1095 <= wire1057[(3'h5):(3'h5)];
              reg1096 <= ({(wire941[(4'hc):(4'hb)] <= ($unsigned(reg1069) ^ wire1056[(3'h4):(3'h4)])),
                      reg1091[(4'he):(1'h0)]} ?
                  (($signed($unsigned(reg1004)) * {(reg1059 ?
                          (7'h48) : reg1093)}) * (^((reg1061 ?
                          reg1008 : reg1077) ?
                      (~reg1015) : $signed(reg1017)))) : reg1092);
            end
          else
            begin
              reg1093 = (+reg1091);
              reg1094 = reg987;
              reg1097 = (8'hb1);
              reg1098 = (wire1055[(3'h6):(3'h4)] ?
                  ($signed($signed({reg1059, wire939})) ^ {(wire942 ?
                          (reg1020 ?
                              (8'hae) : reg1064) : (~&reg1051))}) : $unsigned(forvar1085[(4'h9):(2'h3)]));
            end
        end
      else
        begin
          reg1090 = {(8'hb4)};
          for (forvar1091 = (1'h0); (forvar1091 < (2'h2)); forvar1091 = (forvar1091 + (1'h1)))
            begin
              reg1093 = ($signed(reg1097[(2'h3):(2'h3)]) ?
                  $unsigned($unsigned(reg1074[(3'h7):(3'h5)])) : (&$unsigned($unsigned({(8'ha7),
                      reg1084}))));
              reg1095 <= $signed(((reg982 ?
                      reg1065[(4'ha):(2'h3)] : $unsigned((^reg1086))) ?
                  (~{reg956[(4'he):(4'he)],
                      wire1056[(1'h1):(1'h1)]}) : (reg1092[(3'h4):(1'h0)] >> $signed($signed(reg969)))));
              reg1096 <= wire1056;
              reg1099 <= ((8'ha0) + reg1080);
              reg1100 = $signed(wire938);
            end
          for (forvar1101 = (1'h0); (forvar1101 < (2'h2)); forvar1101 = (forvar1101 + (1'h1)))
            begin
              reg1102 <= reg1070;
              reg1103 = (&((wire1055 >> (+$signed(reg1038))) ^ (reg1013 ?
                  reg956 : (7'h45))));
              reg1104 <= (reg1003 ?
                  $signed((-reg1082[(2'h2):(2'h2)])) : wire1021);
              reg1105 = {((7'h42) < reg1087)};
              reg1106 <= (!reg1104[(5'h11):(1'h0)]);
            end
        end
      reg1107 <= (((~&((reg1074 ?
          forvar1091 : reg1013) || reg1011[(4'h8):(1'h0)])) + $unsigned($signed($unsigned(reg1071)))) == ((~&(^$unsigned(reg1030))) ?
          ((8'ha4) ?
              $signed((reg945 || (7'h46))) : ((reg1087 ? (7'h49) : (7'h48)) ?
                  (reg1008 == reg964) : (!wire940))) : $signed(wire1058[(2'h3):(2'h3)])));
    end
  assign wire1108 = reg969;
  always
    @(posedge clk) begin
      for (forvar1109 = (1'h0); (forvar1109 < (1'h1)); forvar1109 = (forvar1109 + (1'h1)))
        begin
          reg1110 <= $signed($unsigned(reg1026[(3'h5):(2'h3)]));
        end
      for (forvar1111 = (1'h0); (forvar1111 < (2'h2)); forvar1111 = (forvar1111 + (1'h1)))
        begin
          reg1112 <= reg990[(3'h6):(2'h2)];
        end
      reg1113 = ($signed((!((reg1008 ? reg1067 : reg1087) ?
          (reg974 * reg1000) : reg990[(5'h18):(1'h0)]))) == $signed($unsigned(reg1063[(5'h12):(5'h12)])));
      for (forvar1114 = (1'h0); (forvar1114 < (1'h1)); forvar1114 = (forvar1114 + (1'h1)))
        begin
          reg1115 = reg954[(1'h1):(1'h0)];
          reg1116 = (reg955[(2'h2):(2'h2)] ?
              $unsigned(reg1020) : {(($signed(reg1106) | $signed(reg1010)) ^~ {{(7'h49),
                          reg945}})});
          reg1117 <= (($unsigned($unsigned(reg1063[(5'h12):(4'h9)])) ?
              $unsigned((reg1067[(2'h2):(1'h1)] ?
                  reg1030 : $unsigned((8'hbb)))) : $unsigned(((8'h9e) ?
                  $signed(wire1056) : reg1013[(3'h7):(3'h4)]))) >= {(((-reg1026) ?
                  $signed(reg980) : $unsigned((8'ha6))) * $unsigned((reg996 ?
                  reg1049 : wire1060))),
              reg1113[(1'h1):(1'h0)]});
          reg1118 = ((reg1081[(2'h2):(1'h1)] ?
                  $unsigned(wire1108[(4'h8):(3'h7)]) : wire1060[(1'h0):(1'h0)]) ?
              $signed(reg1112) : ($unsigned(reg1000) * $signed(reg1051)));
          for (forvar1119 = (1'h0); (forvar1119 < (3'h4)); forvar1119 = (forvar1119 + (1'h1)))
            begin
              reg1120 <= $signed((7'h40));
              reg1121 <= $signed((+{(~|wire942),
                  {(reg977 ^ forvar1119), (reg1003 ? reg1059 : reg1079)}}));
              reg1122 <= ($signed((~^reg1015[(3'h7):(2'h3)])) >> reg1113[(1'h1):(1'h0)]);
            end
        end
      for (forvar1123 = (1'h0); (forvar1123 < (2'h2)); forvar1123 = (forvar1123 + (1'h1)))
        begin
          reg1124 = reg1095;
          for (forvar1125 = (1'h0); (forvar1125 < (1'h1)); forvar1125 = (forvar1125 + (1'h1)))
            begin
              reg1126 <= (($unsigned((&reg964)) ?
                  (((reg966 <= reg1053) ?
                      (reg961 | wire1060) : reg954[(1'h0):(1'h0)]) < $signed((reg1069 ?
                      (8'haa) : (7'h43)))) : $unsigned((|(wire1056 ?
                      (8'hae) : reg946)))) ~^ $unsigned($unsigned($unsigned(((8'ha1) ?
                  reg1096 : (7'h40))))));
            end
          reg1127 = reg998[(4'h9):(3'h7)];
        end
    end
  always
    @(posedge clk) begin
      reg1128 = $signed(((reg1059[(4'ha):(2'h2)] >= (8'hb8)) >>> (&($signed(reg1088) <= $signed(reg1013)))));
    end
  assign wire1129 = (~reg959[(1'h0):(1'h0)]);
  assign wire1130 = $signed((reg1040 | reg961[(4'hb):(3'h7)]));
  assign wire1131 = ({{(reg1037 ^ (8'ha8))}} ?
                        $signed(($unsigned((reg1038 ? (8'hb2) : reg1003)) ?
                            (-wire939) : reg1030[(1'h1):(1'h0)])) : ($unsigned($signed(reg969)) << $unsigned(reg1078[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      reg1132 <= (|reg996[(3'h5):(1'h0)]);
      for (forvar1133 = (1'h0); (forvar1133 < (2'h2)); forvar1133 = (forvar1133 + (1'h1)))
        begin
          reg1134 <= $unsigned($signed($signed($unsigned(reg1008[(4'h8):(1'h1)]))));
          reg1135 = (+(8'h9c));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module778
#(parameter param871 = ((^~(^~(((8'ha1) ? (8'hbb) : (8'hb0)) ? {(8'h9f), (8'hb1)} : ((8'hb2) >>> (8'haa))))) <= (({(^~(8'hb8)), (^(7'h48))} ^ (+((8'h9e) ? (7'h4a) : (8'h9e)))) >>> (-((|(8'hac)) ? ((7'h4a) ^ (8'haa)) : ((7'h44) != (8'hac)))))))
(y, clk, wire783, wire782, wire781, wire780, wire779);
  output wire [(32'h4d3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire783;
  input wire signed [(5'h12):(1'h0)] wire782;
  input wire [(5'h13):(1'h0)] wire781;
  input wire signed [(3'h7):(1'h0)] wire780;
  input wire [(4'ha):(1'h0)] wire779;
  wire signed [(2'h3):(1'h0)] wire818;
  wire [(2'h2):(1'h0)] wire817;
  wire signed [(5'h17):(1'h0)] wire816;
  reg [(4'he):(1'h0)] reg870 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg869 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg868 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg866 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg864 = (1'h0);
  reg [(5'h11):(1'h0)] reg863 = (1'h0);
  reg [(5'h17):(1'h0)] reg862 = (1'h0);
  reg [(5'h13):(1'h0)] reg858 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg857 = (1'h0);
  reg signed [(4'he):(1'h0)] reg852 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg849 = (1'h0);
  reg [(2'h2):(1'h0)] reg845 = (1'h0);
  reg [(3'h6):(1'h0)] reg838 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg835 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg827 = (1'h0);
  reg [(3'h7):(1'h0)] reg825 = (1'h0);
  reg [(5'h10):(1'h0)] reg822 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg821 = (1'h0);
  reg [(5'h12):(1'h0)] reg820 = (1'h0);
  reg [(3'h7):(1'h0)] reg819 = (1'h0);
  reg [(4'ha):(1'h0)] reg814 = (1'h0);
  reg [(5'h15):(1'h0)] reg813 = (1'h0);
  reg [(4'he):(1'h0)] reg809 = (1'h0);
  reg [(3'h4):(1'h0)] reg807 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg806 = (1'h0);
  reg [(5'h14):(1'h0)] reg804 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg803 = (1'h0);
  reg [(5'h12):(1'h0)] reg802 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg800 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg797 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg796 = (1'h0);
  reg [(3'h4):(1'h0)] reg793 = (1'h0);
  reg [(3'h7):(1'h0)] reg792 = (1'h0);
  reg [(4'ha):(1'h0)] reg790 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg787 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg784 = (1'h0);
  reg [(4'hb):(1'h0)] reg867 = (1'h0);
  reg [(4'h9):(1'h0)] reg865 = (1'h0);
  reg [(3'h5):(1'h0)] forvar863 = (1'h0);
  reg [(5'h16):(1'h0)] reg861 = (1'h0);
  reg [(4'hd):(1'h0)] reg860 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar859 = (1'h0);
  reg [(5'h12):(1'h0)] reg856 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg855 = (1'h0);
  reg [(5'h18):(1'h0)] reg854 = (1'h0);
  reg [(5'h15):(1'h0)] forvar853 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar851 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg850 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg848 = (1'h0);
  reg [(4'hd):(1'h0)] reg847 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg846 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar844 = (1'h0);
  reg [(3'h4):(1'h0)] reg843 = (1'h0);
  reg [(4'hf):(1'h0)] forvar842 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg841 = (1'h0);
  reg [(5'h18):(1'h0)] reg840 = (1'h0);
  reg [(5'h18):(1'h0)] reg839 = (1'h0);
  reg [(4'hb):(1'h0)] reg837 = (1'h0);
  reg [(4'hb):(1'h0)] reg836 = (1'h0);
  reg [(5'h14):(1'h0)] reg834 = (1'h0);
  reg [(5'h11):(1'h0)] forvar833 = (1'h0);
  reg [(4'hd):(1'h0)] reg832 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg831 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg830 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg829 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg828 = (1'h0);
  reg [(4'hc):(1'h0)] forvar824 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg826 = (1'h0);
  reg [(3'h4):(1'h0)] reg824 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg823 = (1'h0);
  reg signed [(4'he):(1'h0)] reg815 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg812 = (1'h0);
  reg [(4'hc):(1'h0)] forvar811 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg810 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg808 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg805 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg801 = (1'h0);
  reg [(2'h3):(1'h0)] reg799 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg798 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar795 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg795 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg794 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg785 = (1'h0);
  reg [(3'h6):(1'h0)] reg791 = (1'h0);
  reg [(5'h13):(1'h0)] reg789 = (1'h0);
  reg [(4'hf):(1'h0)] reg788 = (1'h0);
  reg [(5'h10):(1'h0)] reg786 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar785 = (1'h0);
  assign y = {wire818,
                 wire817,
                 wire816,
                 reg870,
                 reg869,
                 reg868,
                 reg866,
                 reg864,
                 reg863,
                 reg862,
                 reg858,
                 reg857,
                 reg852,
                 reg849,
                 reg845,
                 reg838,
                 reg835,
                 reg827,
                 reg825,
                 reg822,
                 reg821,
                 reg820,
                 reg819,
                 reg814,
                 reg813,
                 reg809,
                 reg807,
                 reg806,
                 reg804,
                 reg803,
                 reg802,
                 reg800,
                 reg797,
                 reg796,
                 reg793,
                 reg792,
                 reg790,
                 reg787,
                 reg784,
                 reg867,
                 reg865,
                 forvar863,
                 reg861,
                 reg860,
                 forvar859,
                 reg856,
                 reg855,
                 reg854,
                 forvar853,
                 forvar851,
                 reg850,
                 reg848,
                 reg847,
                 reg846,
                 forvar844,
                 reg843,
                 forvar842,
                 reg841,
                 reg840,
                 reg839,
                 reg837,
                 reg836,
                 reg834,
                 forvar833,
                 reg832,
                 reg831,
                 reg830,
                 reg829,
                 reg828,
                 forvar824,
                 reg826,
                 reg824,
                 reg823,
                 reg815,
                 reg812,
                 forvar811,
                 reg810,
                 reg808,
                 reg805,
                 reg801,
                 reg799,
                 reg798,
                 forvar795,
                 reg795,
                 reg794,
                 reg785,
                 reg791,
                 reg789,
                 reg788,
                 reg786,
                 forvar785,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ((+{wire781[(4'hc):(4'ha)],
          ({wire779[(2'h3):(1'h0)], {(8'hae), (8'hb6)}} | wire783)}))
        begin
          reg784 <= (wire782[(5'h12):(3'h7)] >>> (wire782[(5'h10):(4'hd)] <= $signed($signed({wire779}))));
          for (forvar785 = (1'h0); (forvar785 < (2'h2)); forvar785 = (forvar785 + (1'h1)))
            begin
              reg786 = (((wire780[(3'h5):(2'h2)] | wire780) ?
                  $signed((wire781[(4'hd):(4'h8)] ?
                      (reg784 ? reg784 : wire779) : (wire780 ?
                          wire779 : forvar785))) : {wire782,
                      $unsigned(wire783[(4'hf):(4'ha)])}) && $signed(((^wire783) ?
                  $unsigned((~&(8'haa))) : $unsigned($unsigned(wire783)))));
              reg787 <= $signed((~&{((wire780 * wire779) ?
                      ((8'hac) & wire779) : (7'h40)),
                  wire782}));
              reg788 = reg786;
              reg789 = reg788[(4'h9):(1'h0)];
              reg790 <= wire782[(4'hc):(3'h5)];
            end
          reg791 = reg788;
        end
      else
        begin
          reg785 = (^~((~^($signed(wire780) ?
              $signed(wire780) : wire782[(4'ha):(4'h9)])) ^ $unsigned($unsigned($signed((8'hb1))))));
          if ((+reg785))
            begin
              reg786 = (-reg785[(3'h7):(3'h4)]);
              reg788 = wire782;
              reg789 = wire782[(3'h4):(2'h2)];
              reg791 = reg787;
            end
          else
            begin
              reg787 <= ($signed(($unsigned($signed(reg790)) ?
                      reg785 : (+(reg786 + wire780)))) ?
                  reg788 : (&{$signed((wire783 ? wire782 : wire783))}));
            end
          reg792 <= reg784;
          reg793 <= {reg785[(2'h3):(1'h0)]};
          reg794 = $signed($signed(($signed($signed(reg792)) ?
              $signed($signed(forvar785)) : $signed(reg791))));
        end
      if (wire780)
        begin
          reg795 = (~^(($signed(forvar785) ?
              $unsigned((-reg789)) : ((reg789 ? wire783 : (7'h48)) ?
                  reg790 : (wire781 ^ forvar785))) - reg787));
        end
      else
        begin
          for (forvar795 = (1'h0); (forvar795 < (2'h3)); forvar795 = (forvar795 + (1'h1)))
            begin
              reg796 <= (-forvar795[(3'h7):(1'h1)]);
              reg797 <= reg787;
              reg798 = ($signed((~^((forvar785 ?
                      wire782 : (8'hb6)) & {reg793}))) ?
                  reg794[(3'h4):(1'h1)] : forvar785[(4'hf):(1'h1)]);
              reg799 = ($signed({(8'ha2),
                  ({reg797, forvar795} ?
                      reg792 : (reg789 * reg798))}) ^~ $unsigned(((reg784[(2'h2):(2'h2)] ?
                  wire781 : reg793[(3'h4):(2'h3)]) >>> ($unsigned(reg797) ?
                  reg796 : ((8'hb8) ? wire780 : wire782)))));
              reg800 <= (8'hb5);
            end
          if (reg794)
            begin
              reg801 = ({(($signed((8'ha0)) >= {reg788,
                          reg795}) && forvar795[(5'h10):(4'hf)]),
                      (reg785[(2'h2):(2'h2)] >>> forvar785)} ?
                  (~(wire782[(2'h3):(1'h1)] | {(-reg795)})) : $signed((((reg788 ?
                      reg791 : reg786) ^~ reg792[(3'h5):(3'h4)]) >> reg797)));
              reg802 <= wire781[(4'hd):(4'hd)];
              reg803 <= wire781[(3'h6):(1'h1)];
              reg804 <= (~&(-forvar785[(4'h8):(1'h0)]));
            end
          else
            begin
              reg801 = $unsigned($signed((reg798[(3'h6):(1'h0)] - reg791)));
              reg805 = ($unsigned(reg802[(4'hb):(4'hb)]) ?
                  (((|reg802[(4'ha):(2'h3)]) ?
                      $unsigned(reg800[(3'h4):(3'h4)]) : (|$signed(wire782))) + $unsigned($unsigned((reg802 | forvar795)))) : $signed(reg793));
              reg806 <= (^~{$unsigned((~&(wire783 & reg796))),
                  $unsigned(((+wire779) ?
                      $signed((7'h40)) : $unsigned(reg794)))});
              reg807 <= {($unsigned($signed((~&reg788))) ^ $signed((reg800[(4'h9):(3'h7)] + $signed(reg791))))};
            end
          reg808 = reg797;
        end
      reg809 <= wire780;
    end
  always
    @(posedge clk) begin
      reg810 = (($signed(wire781) ?
              $unsigned($unsigned({wire783, reg806})) : reg797) ?
          wire779[(3'h5):(2'h2)] : {$unsigned((reg796[(3'h4):(3'h4)] ^ reg792[(3'h7):(3'h7)])),
              ($unsigned((reg787 ? wire779 : reg784)) ^ (!(&wire783)))});
      for (forvar811 = (1'h0); (forvar811 < (2'h2)); forvar811 = (forvar811 + (1'h1)))
        begin
          reg812 = reg784;
          reg813 <= reg804[(3'h5):(2'h3)];
        end
    end
  always
    @(posedge clk) begin
      reg814 <= reg806[(3'h6):(3'h5)];
      reg815 = reg802;
    end
  assign wire816 = (~&($unsigned(($unsigned(reg807) >>> $signed(reg803))) ?
                       $signed($unsigned(reg784[(4'h8):(1'h0)])) : (+$unsigned($unsigned(wire781)))));
  assign wire817 = (wire783 ?
                       (reg797[(1'h1):(1'h0)] & ($unsigned(reg790) != $signed(reg784))) : (reg807 == (reg793[(3'h4):(1'h1)] ?
                           $signed(reg806[(1'h1):(1'h0)]) : (((8'ha9) ?
                                   reg793 : reg813) ?
                               (wire782 ?
                                   reg787 : (8'hb0)) : $signed(reg809)))));
  assign wire818 = reg803[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      if (reg813)
        begin
          if (reg796)
            begin
              reg819 <= ({(^~reg806),
                      {wire780, $unsigned((reg784 == reg806))}} ?
                  {reg806[(3'h4):(2'h2)],
                      ($signed(reg803[(4'hb):(2'h2)]) ?
                          reg803 : reg784)} : $signed(reg804));
              reg820 <= (~^$signed((8'ha2)));
            end
          else
            begin
              reg819 <= (&reg796);
              reg820 <= $unsigned(wire818);
              reg821 <= reg807;
            end
          if ($signed($unsigned(wire783[(4'hc):(2'h2)])))
            begin
              reg822 <= ({$signed(reg796)} >>> ($unsigned($unsigned($unsigned(reg787))) > ($signed((reg819 ?
                      reg814 : reg797)) ?
                  reg807[(1'h1):(1'h0)] : $signed(wire779))));
              reg823 = (wire781 * $signed(reg821[(3'h4):(2'h3)]));
              reg824 = reg822;
              reg825 <= reg822;
            end
          else
            begin
              reg822 <= $unsigned(wire818);
              reg823 = $signed((!wire782[(3'h4):(3'h4)]));
              reg824 = (+(-$signed(reg809[(3'h4):(1'h0)])));
              reg826 = $signed($unsigned((~&{(8'hb2)})));
            end
          reg827 <= (!{$signed(reg793[(1'h1):(1'h0)])});
        end
      else
        begin
          reg823 = reg792[(3'h5):(2'h2)];
          for (forvar824 = (1'h0); (forvar824 < (1'h0)); forvar824 = (forvar824 + (1'h1)))
            begin
              reg826 = {reg797};
              reg828 = (|(8'ha0));
              reg829 = reg813[(5'h13):(4'hc)];
              reg830 = (reg819 ?
                  reg804[(4'he):(3'h4)] : (~$signed($unsigned((~&reg787)))));
            end
        end
      reg831 = ((+$unsigned((-$signed(reg827)))) ?
          (~^reg830) : ((reg822[(4'hf):(3'h7)] || $unsigned($signed(reg822))) ^~ (reg802 ^~ ((~reg809) ?
              $unsigned(reg826) : $unsigned(reg821)))));
      reg832 = reg803;
      for (forvar833 = (1'h0); (forvar833 < (2'h2)); forvar833 = (forvar833 + (1'h1)))
        begin
          if ({$signed(reg797[(1'h1):(1'h1)])})
            begin
              reg834 = {wire816};
              reg835 <= reg803[(3'h4):(1'h0)];
              reg836 = $unsigned({reg813[(5'h15):(4'ha)],
                  (({reg819} ? wire781 : reg807) ?
                      (^~reg832) : (+(wire782 ~^ reg813)))});
            end
          else
            begin
              reg834 = reg824;
              reg836 = $signed(wire779);
              reg837 = reg824;
              reg838 <= $signed(wire782[(3'h7):(3'h7)]);
            end
          if ($signed($signed(wire780[(3'h7):(1'h0)])))
            begin
              reg839 = $signed($unsigned($signed(((~&reg829) ?
                  (reg837 ^ reg802) : reg829[(4'ha):(3'h5)]))));
            end
          else
            begin
              reg839 = reg784[(2'h3):(2'h3)];
              reg840 = $signed(reg822);
            end
          reg841 = $unsigned($unsigned(reg784));
        end
      for (forvar842 = (1'h0); (forvar842 < (3'h4)); forvar842 = (forvar842 + (1'h1)))
        begin
          reg843 = (^$unsigned(({reg792} == (^$unsigned(reg834)))));
          for (forvar844 = (1'h0); (forvar844 < (2'h2)); forvar844 = (forvar844 + (1'h1)))
            begin
              reg845 <= (~^$signed(wire779));
              reg846 = reg809;
              reg847 = $signed($unsigned((reg819[(3'h6):(3'h5)] ?
                  $unsigned($signed(reg843)) : {$signed(reg792), reg784})));
              reg848 = ($unsigned($signed(reg784[(2'h2):(1'h0)])) >= (|reg837));
            end
          reg849 <= $signed((&(8'hb2)));
        end
    end
  always
    @(posedge clk) begin
      reg850 = (8'hae);
      for (forvar851 = (1'h0); (forvar851 < (2'h3)); forvar851 = (forvar851 + (1'h1)))
        begin
          reg852 <= ({$signed((+(reg835 ~^ reg796))), reg820[(4'h8):(4'h8)]} ?
              $signed(reg787[(3'h7):(3'h6)]) : reg797);
          for (forvar853 = (1'h0); (forvar853 < (1'h0)); forvar853 = (forvar853 + (1'h1)))
            begin
              reg854 = $signed(reg825[(3'h6):(2'h3)]);
              reg855 = reg797[(1'h0):(1'h0)];
              reg856 = ((&{$signed((reg802 ? reg825 : reg821))}) ?
                  $signed((|forvar851)) : reg802);
              reg857 <= reg814[(2'h2):(1'h1)];
            end
          reg858 <= (~$signed((^reg857[(4'h8):(2'h2)])));
          for (forvar859 = (1'h0); (forvar859 < (3'h4)); forvar859 = (forvar859 + (1'h1)))
            begin
              reg860 = reg813[(3'h5):(3'h5)];
              reg861 = (~{(((reg852 >>> reg813) ?
                          $signed((7'h43)) : $unsigned(reg838)) ?
                      $signed($signed(reg804)) : ($signed(forvar859) ?
                          reg827[(2'h2):(1'h0)] : $unsigned((7'h46))))});
            end
        end
      reg862 <= ($signed((&(reg838 ?
          reg857[(1'h0):(1'h0)] : ((8'ha1) ?
              reg804 : (8'hae))))) ^~ $signed(($signed($signed(wire782)) + ($unsigned(forvar859) ?
          reg857[(1'h0):(1'h0)] : ((8'ha7) ? reg849 : reg790)))));
      if ($signed(({(7'h42), reg803[(3'h5):(3'h4)]} ?
          {(!(reg792 ? (8'hb9) : (8'hb9))),
              {(reg861 ? (8'ha6) : (8'hac))}} : ((^~wire818[(2'h3):(2'h3)]) ?
              $signed($signed(forvar859)) : ($signed((8'ha6)) ?
                  forvar859[(4'he):(3'h4)] : (reg784 || (7'h4a)))))))
        begin
          reg863 <= $unsigned(reg856[(3'h7):(3'h5)]);
        end
      else
        begin
          for (forvar863 = (1'h0); (forvar863 < (1'h0)); forvar863 = (forvar863 + (1'h1)))
            begin
              reg864 <= (reg845[(1'h1):(1'h1)] ?
                  reg809[(4'ha):(2'h2)] : (^~(~^wire783)));
            end
          if (($signed(reg863) ?
              ((($unsigned(reg849) ~^ (~^reg809)) ?
                      $signed(reg852[(3'h7):(3'h4)]) : forvar863[(1'h1):(1'h1)]) ?
                  {((!reg819) ?
                          {(8'hbc), wire816} : (reg856 ?
                              reg838 : (7'h48)))} : forvar859[(4'h9):(4'h9)]) : forvar851[(1'h0):(1'h0)]))
            begin
              reg865 = reg797[(2'h3):(1'h0)];
              reg866 <= wire816;
              reg867 = (~|(^$unsigned(reg822)));
            end
          else
            begin
              reg866 <= (!wire779);
              reg868 <= $unsigned(($unsigned(reg807[(1'h0):(1'h0)]) >>> reg827[(3'h4):(3'h4)]));
              reg869 <= (($unsigned((((8'hbb) >>> reg849) ^~ {(8'hbf)})) ?
                  reg850[(4'hf):(4'h8)] : $signed(($unsigned(reg797) <= $signed((8'hb0))))) >= ({(~|{forvar859})} * ($unsigned((reg792 ?
                      reg792 : (8'ha7))) ?
                  reg784 : $unsigned($unsigned((7'h45))))));
            end
          reg870 <= ((~|(((reg854 + forvar853) - reg835) ?
                  (&reg866) : {$signed((8'hb4)), reg807})) ?
              (7'h43) : $unsigned($signed(reg806)));
        end
    end
endmodule