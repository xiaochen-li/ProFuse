(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'hfa9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire3;
  input wire [(5'h15):(1'h0)] wire2;
  input wire [(5'h17):(1'h0)] wire1;
  input wire signed [(4'hc):(1'h0)] wire0;
  wire signed [(4'ha):(1'h0)] wire1492;
  wire signed [(5'h17):(1'h0)] wire1467;
  wire [(5'h11):(1'h0)] wire272;
  wire [(4'he):(1'h0)] wire271;
  wire signed [(5'h14):(1'h0)] wire270;
  wire signed [(2'h3):(1'h0)] wire190;
  wire [(3'h6):(1'h0)] wire189;
  wire signed [(5'h18):(1'h0)] wire188;
  wire signed [(5'h17):(1'h0)] wire186;
  wire signed [(5'h12):(1'h0)] wire185;
  wire [(5'h13):(1'h0)] wire184;
  wire [(4'hc):(1'h0)] wire63;
  wire signed [(5'h11):(1'h0)] wire4;
  reg [(5'h16):(1'h0)] reg1489 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1488 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1487 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1485 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1484 = (1'h0);
  reg [(5'h12):(1'h0)] reg1481 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1480 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1479 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1475 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1473 = (1'h0);
  reg [(3'h7):(1'h0)] reg1472 = (1'h0);
  reg [(4'ha):(1'h0)] reg1471 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg7 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg10 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg11 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg13 = (1'h0);
  reg [(4'h9):(1'h0)] reg15 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg16 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg17 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg22 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg6 = (1'h0);
  reg [(3'h4):(1'h0)] reg23 = (1'h0);
  reg [(2'h2):(1'h0)] reg26 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg29 = (1'h0);
  reg [(5'h18):(1'h0)] reg30 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg32 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg37 = (1'h0);
  reg [(4'hf):(1'h0)] reg38 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg39 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg41 = (1'h0);
  reg [(5'h12):(1'h0)] reg43 = (1'h0);
  reg [(5'h14):(1'h0)] reg44 = (1'h0);
  reg [(5'h11):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg50 = (1'h0);
  reg [(4'he):(1'h0)] reg52 = (1'h0);
  reg [(5'h11):(1'h0)] reg53 = (1'h0);
  reg [(5'h12):(1'h0)] reg55 = (1'h0);
  reg [(5'h12):(1'h0)] reg56 = (1'h0);
  reg [(5'h15):(1'h0)] reg58 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg60 = (1'h0);
  reg [(5'h14):(1'h0)] reg61 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg62 = (1'h0);
  reg signed [(4'he):(1'h0)] reg64 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg70 = (1'h0);
  reg [(4'h9):(1'h0)] reg72 = (1'h0);
  reg [(5'h16):(1'h0)] reg74 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg75 = (1'h0);
  reg [(5'h17):(1'h0)] reg77 = (1'h0);
  reg [(4'hf):(1'h0)] reg78 = (1'h0);
  reg [(5'h16):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg87 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg89 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg92 = (1'h0);
  reg [(5'h16):(1'h0)] reg97 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg100 = (1'h0);
  reg [(4'h8):(1'h0)] reg102 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg105 = (1'h0);
  reg [(3'h4):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg110 = (1'h0);
  reg [(5'h13):(1'h0)] reg113 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg115 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg116 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg117 = (1'h0);
  reg [(4'hf):(1'h0)] reg119 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg122 = (1'h0);
  reg [(4'h8):(1'h0)] reg125 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg126 = (1'h0);
  reg [(5'h10):(1'h0)] reg130 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg133 = (1'h0);
  reg [(4'hc):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg136 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg139 = (1'h0);
  reg [(4'hb):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg148 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg150 = (1'h0);
  reg [(2'h3):(1'h0)] reg152 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg154 = (1'h0);
  reg signed [(4'he):(1'h0)] reg156 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg157 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg158 = (1'h0);
  reg [(5'h13):(1'h0)] reg159 = (1'h0);
  reg [(2'h3):(1'h0)] reg163 = (1'h0);
  reg [(5'h13):(1'h0)] reg165 = (1'h0);
  reg [(3'h4):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg170 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg172 = (1'h0);
  reg [(3'h4):(1'h0)] reg175 = (1'h0);
  reg [(4'hd):(1'h0)] reg177 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg179 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg181 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg183 = (1'h0);
  reg [(5'h17):(1'h0)] reg187 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg193 = (1'h0);
  reg [(3'h5):(1'h0)] reg194 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg195 = (1'h0);
  reg [(4'ha):(1'h0)] reg196 = (1'h0);
  reg [(2'h3):(1'h0)] reg197 = (1'h0);
  reg [(3'h7):(1'h0)] reg199 = (1'h0);
  reg [(4'h8):(1'h0)] reg201 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg202 = (1'h0);
  reg signed [(4'he):(1'h0)] reg203 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg205 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg206 = (1'h0);
  reg [(4'he):(1'h0)] reg208 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg212 = (1'h0);
  reg [(3'h5):(1'h0)] reg214 = (1'h0);
  reg [(5'h16):(1'h0)] reg215 = (1'h0);
  reg [(4'hd):(1'h0)] reg217 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg220 = (1'h0);
  reg [(4'hf):(1'h0)] reg223 = (1'h0);
  reg [(5'h11):(1'h0)] reg228 = (1'h0);
  reg signed [(4'he):(1'h0)] reg229 = (1'h0);
  reg [(2'h3):(1'h0)] reg231 = (1'h0);
  reg [(4'h9):(1'h0)] reg235 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg241 = (1'h0);
  reg [(4'ha):(1'h0)] reg246 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg247 = (1'h0);
  reg [(5'h10):(1'h0)] reg248 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg255 = (1'h0);
  reg signed [(4'he):(1'h0)] reg258 = (1'h0);
  reg [(5'h10):(1'h0)] reg260 = (1'h0);
  reg [(5'h13):(1'h0)] reg262 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg268 = (1'h0);
  reg [(4'he):(1'h0)] reg1491 = (1'h0);
  reg [(3'h7):(1'h0)] reg1490 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1486 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1483 = (1'h0);
  reg [(3'h6):(1'h0)] reg1482 = (1'h0);
  reg [(4'h9):(1'h0)] reg1478 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1477 = (1'h0);
  reg [(4'hd):(1'h0)] reg1476 = (1'h0);
  reg [(5'h16):(1'h0)] reg1474 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1470 = (1'h0);
  reg [(4'hb):(1'h0)] reg1469 = (1'h0);
  reg [(4'hc):(1'h0)] reg269 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar267 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg266 = (1'h0);
  reg [(2'h2):(1'h0)] reg265 = (1'h0);
  reg [(4'h9):(1'h0)] forvar264 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg263 = (1'h0);
  reg [(4'hc):(1'h0)] forvar257 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg261 = (1'h0);
  reg [(5'h18):(1'h0)] reg259 = (1'h0);
  reg [(4'hc):(1'h0)] reg257 = (1'h0);
  reg [(4'hf):(1'h0)] reg256 = (1'h0);
  reg [(5'h14):(1'h0)] reg254 = (1'h0);
  reg [(4'hd):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg252 = (1'h0);
  reg [(2'h3):(1'h0)] reg251 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg250 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg245 = (1'h0);
  reg [(3'h5):(1'h0)] reg244 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg243 = (1'h0);
  reg [(4'hf):(1'h0)] reg242 = (1'h0);
  reg [(3'h6):(1'h0)] forvar239 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg238 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar237 = (1'h0);
  reg [(5'h17):(1'h0)] reg236 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg234 = (1'h0);
  reg [(3'h7):(1'h0)] reg233 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar232 = (1'h0);
  reg signed [(4'he):(1'h0)] reg230 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar227 = (1'h0);
  reg [(4'hf):(1'h0)] reg226 = (1'h0);
  reg [(5'h10):(1'h0)] reg225 = (1'h0);
  reg [(2'h3):(1'h0)] reg224 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg222 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar221 = (1'h0);
  reg [(4'hb):(1'h0)] reg219 = (1'h0);
  reg [(4'he):(1'h0)] forvar218 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar216 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar213 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg211 = (1'h0);
  reg [(4'h8):(1'h0)] reg210 = (1'h0);
  reg signed [(4'he):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar207 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg200 = (1'h0);
  reg [(4'he):(1'h0)] forvar194 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar200 = (1'h0);
  reg [(2'h3):(1'h0)] reg198 = (1'h0);
  reg [(5'h12):(1'h0)] reg192 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg191 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg180 = (1'h0);
  reg [(5'h11):(1'h0)] forvar178 = (1'h0);
  reg [(5'h15):(1'h0)] reg176 = (1'h0);
  reg [(2'h2):(1'h0)] reg174 = (1'h0);
  reg [(5'h10):(1'h0)] reg173 = (1'h0);
  reg [(5'h10):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg169 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg168 = (1'h0);
  reg [(4'hb):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar164 = (1'h0);
  reg [(4'ha):(1'h0)] reg162 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg161 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg160 = (1'h0);
  reg [(4'hf):(1'h0)] reg155 = (1'h0);
  reg signed [(4'he):(1'h0)] reg153 = (1'h0);
  reg [(5'h16):(1'h0)] forvar151 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg149 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar146 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg144 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar143 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg142 = (1'h0);
  reg [(3'h6):(1'h0)] reg141 = (1'h0);
  reg [(5'h18):(1'h0)] reg140 = (1'h0);
  reg [(4'ha):(1'h0)] reg138 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg137 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg135 = (1'h0);
  reg [(5'h18):(1'h0)] reg132 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg131 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg129 = (1'h0);
  reg [(5'h18):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg127 = (1'h0);
  reg [(4'he):(1'h0)] reg124 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg123 = (1'h0);
  reg [(5'h15):(1'h0)] forvar119 = (1'h0);
  reg [(3'h7):(1'h0)] reg112 = (1'h0);
  reg [(5'h13):(1'h0)] forvar111 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg121 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg120 = (1'h0);
  reg [(4'hd):(1'h0)] reg118 = (1'h0);
  reg [(2'h2):(1'h0)] reg114 = (1'h0);
  reg [(4'he):(1'h0)] forvar112 = (1'h0);
  reg [(4'ha):(1'h0)] reg111 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg108 = (1'h0);
  reg [(5'h12):(1'h0)] forvar106 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar102 = (1'h0);
  reg [(5'h14):(1'h0)] reg104 = (1'h0);
  reg [(4'h8):(1'h0)] reg103 = (1'h0);
  reg [(5'h10):(1'h0)] reg101 = (1'h0);
  reg [(4'hb):(1'h0)] reg99 = (1'h0);
  reg [(3'h7):(1'h0)] reg98 = (1'h0);
  reg [(4'hd):(1'h0)] reg96 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg95 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg94 = (1'h0);
  reg [(3'h7):(1'h0)] reg93 = (1'h0);
  reg [(3'h4):(1'h0)] reg91 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar90 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg86 = (1'h0);
  reg [(5'h14):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar84 = (1'h0);
  reg [(2'h2):(1'h0)] reg83 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg82 = (1'h0);
  reg [(5'h13):(1'h0)] forvar81 = (1'h0);
  reg [(4'ha):(1'h0)] reg80 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg73 = (1'h0);
  reg [(5'h10):(1'h0)] reg71 = (1'h0);
  reg [(4'he):(1'h0)] reg68 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg66 = (1'h0);
  reg [(5'h15):(1'h0)] reg65 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg59 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar57 = (1'h0);
  reg [(5'h15):(1'h0)] reg54 = (1'h0);
  reg [(4'ha):(1'h0)] reg51 = (1'h0);
  reg [(2'h3):(1'h0)] forvar49 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg48 = (1'h0);
  reg [(3'h7):(1'h0)] forvar47 = (1'h0);
  reg [(4'hc):(1'h0)] reg46 = (1'h0);
  reg [(3'h4):(1'h0)] reg42 = (1'h0);
  reg [(5'h15):(1'h0)] forvar38 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar28 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar23 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg40 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg36 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg35 = (1'h0);
  reg [(4'hc):(1'h0)] reg34 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg33 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg31 = (1'h0);
  reg [(4'hb):(1'h0)] reg28 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg27 = (1'h0);
  reg [(4'h9):(1'h0)] reg25 = (1'h0);
  reg [(2'h3):(1'h0)] reg24 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar14 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar12 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar7 = (1'h0);
  reg [(2'h2):(1'h0)] reg21 = (1'h0);
  reg [(4'h8):(1'h0)] reg20 = (1'h0);
  reg [(5'h11):(1'h0)] reg18 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg14 = (1'h0);
  reg [(5'h16):(1'h0)] reg12 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg9 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg8 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar6 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg5 = (1'h0);
  assign y = {wire1492,
                 wire1467,
                 wire272,
                 wire271,
                 wire270,
                 wire190,
                 wire189,
                 wire188,
                 wire186,
                 wire185,
                 wire184,
                 wire63,
                 wire4,
                 reg1489,
                 reg1488,
                 reg1487,
                 reg1485,
                 reg1484,
                 reg1481,
                 reg1480,
                 reg1479,
                 reg1475,
                 reg1473,
                 reg1472,
                 reg1471,
                 reg7,
                 reg10,
                 reg11,
                 reg13,
                 reg15,
                 reg16,
                 reg17,
                 reg19,
                 reg22,
                 reg6,
                 reg23,
                 reg26,
                 reg29,
                 reg30,
                 reg32,
                 reg37,
                 reg38,
                 reg39,
                 reg41,
                 reg43,
                 reg44,
                 reg45,
                 reg50,
                 reg52,
                 reg53,
                 reg55,
                 reg56,
                 reg58,
                 reg60,
                 reg61,
                 reg62,
                 reg64,
                 reg69,
                 reg70,
                 reg72,
                 reg74,
                 reg75,
                 reg77,
                 reg78,
                 reg79,
                 reg87,
                 reg88,
                 reg89,
                 reg92,
                 reg97,
                 reg100,
                 reg102,
                 reg90,
                 reg105,
                 reg107,
                 reg109,
                 reg110,
                 reg113,
                 reg115,
                 reg116,
                 reg117,
                 reg119,
                 reg122,
                 reg125,
                 reg126,
                 reg130,
                 reg133,
                 reg134,
                 reg136,
                 reg139,
                 reg145,
                 reg148,
                 reg150,
                 reg152,
                 reg154,
                 reg156,
                 reg157,
                 reg158,
                 reg159,
                 reg163,
                 reg165,
                 reg166,
                 reg170,
                 reg172,
                 reg175,
                 reg177,
                 reg179,
                 reg181,
                 reg182,
                 reg183,
                 reg187,
                 reg193,
                 reg194,
                 reg195,
                 reg196,
                 reg197,
                 reg199,
                 reg201,
                 reg202,
                 reg203,
                 reg205,
                 reg206,
                 reg208,
                 reg212,
                 reg214,
                 reg215,
                 reg217,
                 reg220,
                 reg223,
                 reg228,
                 reg229,
                 reg231,
                 reg235,
                 reg240,
                 reg241,
                 reg246,
                 reg247,
                 reg248,
                 reg255,
                 reg258,
                 reg260,
                 reg262,
                 reg268,
                 reg1491,
                 reg1490,
                 reg1486,
                 reg1483,
                 reg1482,
                 reg1478,
                 reg1477,
                 reg1476,
                 reg1474,
                 reg1470,
                 reg1469,
                 reg269,
                 forvar267,
                 reg266,
                 reg265,
                 forvar264,
                 reg263,
                 forvar257,
                 reg261,
                 reg259,
                 reg257,
                 reg256,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 forvar239,
                 reg238,
                 forvar237,
                 reg236,
                 reg234,
                 reg233,
                 forvar232,
                 reg230,
                 forvar227,
                 reg226,
                 reg225,
                 reg224,
                 reg222,
                 forvar221,
                 reg219,
                 forvar218,
                 forvar216,
                 forvar213,
                 reg211,
                 reg210,
                 reg209,
                 forvar207,
                 reg200,
                 forvar194,
                 reg204,
                 forvar200,
                 reg198,
                 reg192,
                 reg191,
                 reg180,
                 forvar178,
                 reg176,
                 reg174,
                 reg173,
                 reg171,
                 reg169,
                 reg168,
                 reg167,
                 forvar164,
                 reg162,
                 reg161,
                 reg160,
                 reg155,
                 reg153,
                 forvar151,
                 reg149,
                 reg147,
                 forvar146,
                 reg144,
                 forvar143,
                 reg142,
                 reg141,
                 reg140,
                 reg138,
                 reg137,
                 reg135,
                 reg132,
                 reg131,
                 reg129,
                 reg128,
                 reg127,
                 reg124,
                 reg123,
                 forvar119,
                 reg112,
                 forvar111,
                 reg121,
                 reg120,
                 reg118,
                 reg114,
                 forvar112,
                 reg111,
                 reg108,
                 forvar106,
                 forvar102,
                 reg104,
                 reg103,
                 reg101,
                 reg99,
                 reg98,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg91,
                 forvar90,
                 reg86,
                 reg85,
                 forvar84,
                 reg83,
                 reg82,
                 forvar81,
                 reg80,
                 reg76,
                 reg73,
                 reg71,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg59,
                 forvar57,
                 reg54,
                 reg51,
                 forvar49,
                 reg48,
                 forvar47,
                 reg46,
                 reg42,
                 forvar38,
                 forvar28,
                 forvar23,
                 reg40,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg31,
                 reg28,
                 reg27,
                 reg25,
                 reg24,
                 forvar14,
                 forvar12,
                 forvar7,
                 reg21,
                 reg20,
                 reg18,
                 reg14,
                 reg12,
                 reg9,
                 reg8,
                 forvar6,
                 reg5,
                 (1'h0)};
  assign wire4 = $signed(((wire0 ? wire1 : (|wire0)) ?
                     (&(~^$unsigned((7'h43)))) : $signed(wire3)));
  always
    @(posedge clk) begin
      if ({wire0[(4'ha):(2'h2)]})
        begin
          reg5 = $unsigned($signed($unsigned($signed($signed(wire2)))));
          for (forvar6 = (1'h0); (forvar6 < (2'h2)); forvar6 = (forvar6 + (1'h1)))
            begin
              reg7 <= ($signed(($unsigned((^~wire4)) > ($signed(forvar6) ?
                      (wire3 != forvar6) : $signed(forvar6)))) ?
                  $unsigned(wire3) : wire2[(1'h1):(1'h1)]);
            end
          if ((wire3[(3'h6):(3'h6)] >= ($signed($signed($signed(wire3))) ?
              $unsigned($unsigned(((8'h9e) << wire4))) : ((((8'hb7) | forvar6) ?
                      (~|wire3) : (wire0 ? (8'hbd) : reg5)) ?
                  (~|$unsigned(wire4)) : ((wire1 > reg5) << reg5[(3'h4):(1'h0)])))))
            begin
              reg8 = $unsigned(($signed(wire4) || $unsigned((~&$signed(wire4)))));
              reg9 = ($signed(({wire4[(1'h0):(1'h0)]} ^~ (-((7'h45) ?
                      wire3 : wire1)))) ?
                  (^wire2[(1'h0):(1'h0)]) : reg5);
            end
          else
            begin
              reg10 <= forvar6;
              reg11 <= (({$signed(wire1),
                          ((reg9 * reg7) ? wire4 : $signed(wire2))} ?
                      $signed(((forvar6 <= wire2) <= $signed(forvar6))) : ({$signed(wire3),
                              (wire3 ? (8'hab) : wire1)} ?
                          {(~wire0)} : $unsigned((-reg10)))) ?
                  $signed((^~reg10[(3'h4):(2'h2)])) : (reg9[(3'h4):(2'h3)] ?
                      $unsigned((-(reg5 >= wire2))) : $unsigned(wire1)));
              reg12 = wire1[(1'h1):(1'h0)];
              reg13 <= $unsigned(reg7);
              reg14 = reg9;
            end
          if ($signed({(-reg14), $unsigned(reg14)}))
            begin
              reg15 <= wire4[(2'h2):(1'h0)];
              reg16 <= reg9[(2'h3):(1'h1)];
              reg17 <= ({{reg11}} >>> ($signed($unsigned((^~(8'h9f)))) >= $signed(reg10[(2'h2):(1'h1)])));
              reg18 = reg14;
              reg19 <= ($signed((7'h40)) ?
                  $signed((((~&reg13) > (wire4 ^~ reg16)) ?
                      $unsigned((&wire3)) : (!reg12))) : reg7);
            end
          else
            begin
              reg18 = wire3[(5'h11):(4'hf)];
              reg19 <= forvar6[(4'hb):(4'h8)];
              reg20 = $unsigned((-forvar6));
              reg21 = wire4[(4'h9):(2'h2)];
              reg22 <= (&reg15);
            end
        end
      else
        begin
          reg5 = (reg14[(2'h2):(1'h0)] * wire0[(3'h7):(3'h5)]);
          reg6 <= reg14[(1'h0):(1'h0)];
          for (forvar7 = (1'h0); (forvar7 < (2'h3)); forvar7 = (forvar7 + (1'h1)))
            begin
              reg10 <= (wire1 ? (~|reg10) : $signed(forvar7));
              reg11 <= ($signed($signed((~&(-forvar7)))) - $unsigned((((reg15 ?
                      reg17 : (8'hb3)) ?
                  (reg15 >= reg18) : $signed(reg18)) > ($signed(reg16) ?
                  $signed(reg18) : (reg18 ? reg19 : (8'hb8))))));
            end
          for (forvar12 = (1'h0); (forvar12 < (1'h0)); forvar12 = (forvar12 + (1'h1)))
            begin
              reg13 <= ($unsigned(reg13) ^ $unsigned(({reg17[(2'h2):(1'h0)]} << (!forvar7))));
            end
          for (forvar14 = (1'h0); (forvar14 < (1'h0)); forvar14 = (forvar14 + (1'h1)))
            begin
              reg15 <= reg11;
              reg16 <= (reg22[(2'h3):(1'h0)] * $signed($unsigned($unsigned((wire3 ?
                  reg21 : (8'hbd))))));
              reg18 = ($unsigned(($signed(reg6) ?
                      $signed($unsigned(reg19)) : forvar6)) ?
                  $signed(reg17[(3'h6):(3'h5)]) : {forvar14,
                      {$signed((!reg11)),
                          $unsigned((reg21 ? forvar6 : forvar6))}});
              reg20 = wire0[(1'h1):(1'h0)];
            end
        end
      if ($signed((({(~^wire3), (~|reg7)} ?
              (|reg17[(2'h3):(1'h1)]) : $signed($signed(wire4))) ?
          reg6[(4'h9):(3'h7)] : (((reg9 ? reg8 : reg5) - $signed((8'haa))) ?
              reg15[(1'h1):(1'h0)] : reg6))))
        begin
          if ($unsigned(reg10))
            begin
              reg23 <= {({$unsigned((wire1 ?
                          wire3 : reg18))} && ((^~reg10[(3'h5):(3'h4)]) ?
                      reg11 : reg20)),
                  reg7[(4'h9):(3'h5)]};
              reg24 = $unsigned({({(7'h48)} ? reg20 : $unsigned((-reg22)))});
            end
          else
            begin
              reg24 = (&$signed(reg24[(1'h0):(1'h0)]));
              reg25 = (!reg21[(1'h1):(1'h1)]);
              reg26 <= reg6;
              reg27 = ((|({$signed(wire0),
                      reg18[(4'hc):(3'h7)]} << $signed((reg6 ?
                      reg13 : reg6)))) ?
                  forvar6 : reg9);
              reg28 = (^~reg22);
            end
          reg29 <= $unsigned($signed($unsigned((((8'haa) + reg27) ^~ (reg16 ?
              reg15 : reg18)))));
          if ($unsigned(reg17[(1'h0):(1'h0)]))
            begin
              reg30 <= reg10;
            end
          else
            begin
              reg31 = {(^(~&({reg11} <= (reg11 ^~ forvar6))))};
              reg32 <= reg23;
              reg33 = (!(($signed(reg30[(5'h14):(3'h6)]) - forvar6) >= (&(reg24 - $unsigned((8'h9d))))));
              reg34 = wire0;
            end
          if ({(&forvar7),
              ((~&$unsigned((reg12 ? reg16 : reg19))) ?
                  {(~|wire3), ((reg22 ^~ reg19) <= {reg33})} : reg7)})
            begin
              reg35 = $signed(((+(wire4[(3'h7):(3'h7)] ?
                      reg15 : reg7[(5'h12):(1'h1)])) ?
                  {reg15,
                      ((^~forvar6) == $unsigned(wire1))} : (($signed(wire3) != reg18) == ($signed((8'h9f)) ?
                      $unsigned(reg5) : $signed(reg30)))));
              reg36 = reg22[(3'h5):(2'h3)];
            end
          else
            begin
              reg37 <= {reg17[(1'h1):(1'h1)],
                  $signed((wire1 ?
                      (^reg23[(2'h3):(2'h2)]) : ({(8'ha8), reg17} ?
                          (reg11 << (8'ha6)) : reg17[(1'h0):(1'h0)])))};
              reg38 <= $unsigned((reg5 == $unsigned((reg32 == (reg20 ?
                  reg23 : wire3)))));
              reg39 <= reg23[(1'h1):(1'h0)];
              reg40 = {$signed($unsigned($unsigned(reg38))), {reg5, reg31}};
              reg41 <= (8'had);
            end
        end
      else
        begin
          for (forvar23 = (1'h0); (forvar23 < (1'h0)); forvar23 = (forvar23 + (1'h1)))
            begin
              reg24 = ((!(((forvar6 || reg19) ?
                          reg6[(4'h9):(4'h9)] : (~&reg30)) ?
                      $unsigned($signed(forvar14)) : ((reg18 ~^ (7'h40)) <= (reg27 ?
                          reg31 : reg15)))) ?
                  ((~|reg40) - (8'ha6)) : (reg35[(5'h11):(4'ha)] << (~$unsigned((&reg16)))));
              reg26 <= reg29[(2'h3):(1'h1)];
              reg27 = (({reg20[(4'h8):(3'h6)]} ?
                  (reg40 ^~ (&wire4[(3'h7):(2'h2)])) : (((reg28 * wire3) >>> (reg13 && (8'hba))) * {(&wire0),
                      reg41})) <<< $signed(reg21[(2'h2):(1'h1)]));
            end
          for (forvar28 = (1'h0); (forvar28 < (2'h2)); forvar28 = (forvar28 + (1'h1)))
            begin
              reg31 = (reg10 ?
                  ($unsigned(((reg17 & (8'hb0)) ?
                          reg5 : reg15[(3'h5):(1'h1)])) ?
                      $signed($unsigned((reg36 & (7'h48)))) : (reg29[(2'h2):(1'h0)] != reg40[(4'hb):(4'h8)])) : {reg26[(1'h1):(1'h1)],
                      reg8[(5'h10):(4'hf)]});
              reg32 <= reg18;
              reg33 = {reg18[(4'hf):(4'hd)], (^$unsigned((~(8'hbf))))};
              reg37 <= reg14[(1'h1):(1'h0)];
            end
          for (forvar38 = (1'h0); (forvar38 < (2'h2)); forvar38 = (forvar38 + (1'h1)))
            begin
              reg39 <= ($unsigned($signed((7'h43))) ?
                  $signed((~^$unsigned((8'hbe)))) : (reg25[(2'h3):(1'h1)] ?
                      (~|(reg33 && reg33)) : $unsigned((|$unsigned((7'h44))))));
              reg41 <= $signed((~&$signed((reg26[(1'h0):(1'h0)] ?
                  (reg7 ? reg7 : reg39) : (~^(8'h9c))))));
              reg42 = forvar14[(2'h2):(1'h1)];
              reg43 <= (reg12 + $unsigned(((reg7 ? (^~wire3) : forvar14) ?
                  ({reg20,
                      (8'hb0)} * $unsigned(reg22)) : $unsigned(reg11[(2'h2):(2'h2)]))));
            end
          reg44 <= $unsigned(($signed($unsigned($unsigned(reg22))) ?
              reg23[(2'h2):(1'h1)] : $unsigned(((reg27 ? reg13 : reg38) ?
                  (wire0 == wire4) : reg14[(2'h2):(1'h0)]))));
          if ($unsigned($signed($signed((~&((8'hb1) | (8'ha3)))))))
            begin
              reg45 <= $unsigned((~&$unsigned(wire3[(3'h6):(1'h0)])));
            end
          else
            begin
              reg46 = forvar6;
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar47 = (1'h0); (forvar47 < (1'h1)); forvar47 = (forvar47 + (1'h1)))
        begin
          reg48 = ($unsigned($signed((~&reg29))) != (reg37[(3'h7):(2'h3)] ^~ (^reg22)));
          for (forvar49 = (1'h0); (forvar49 < (1'h0)); forvar49 = (forvar49 + (1'h1)))
            begin
              reg50 <= reg16;
            end
        end
      if (reg10)
        begin
          reg51 = {(-reg22)};
        end
      else
        begin
          reg51 = $unsigned(wire4[(3'h6):(2'h2)]);
          if (({$signed(reg17[(3'h7):(3'h7)]),
              reg38} && $unsigned($signed(wire0))))
            begin
              reg52 <= $signed(((($signed(reg17) >= $signed((7'h44))) == $signed((reg19 && reg17))) ?
                  (reg26 > $signed($unsigned((7'h49)))) : {reg22[(3'h5):(2'h3)]}));
              reg53 <= ($signed(reg6[(2'h2):(2'h2)]) ?
                  ((&((~^wire3) ?
                      $unsigned(reg45) : $unsigned(reg16))) + {((-(8'ha3)) ?
                          $unsigned(reg29) : $signed(reg10))}) : $signed({{reg17}}));
            end
          else
            begin
              reg52 <= ((reg37[(3'h7):(3'h6)] ?
                      (reg44[(4'hc):(1'h1)] >= $signed($signed(wire3))) : reg53[(3'h7):(3'h5)]) ?
                  (reg38[(4'hd):(3'h7)] <<< ((|reg15[(3'h4):(1'h0)]) >= $unsigned(reg32))) : {$unsigned($signed(((8'hb1) < (7'h40))))});
              reg53 <= (reg16 <<< reg48[(1'h1):(1'h0)]);
              reg54 = (({(+$signed(reg11))} ^ {wire1}) >>> (-(^((reg13 ?
                  reg37 : reg15) >> reg30))));
              reg55 <= $signed($signed((((reg29 ? reg13 : wire4) ?
                  reg51[(1'h1):(1'h0)] : (|wire3)) != $unsigned($unsigned(reg11)))));
              reg56 <= (((({(7'h45)} > (!(8'hbf))) ?
                  {$signed(reg54)} : ((wire1 ? reg44 : wire3) ?
                      wire4[(3'h7):(1'h0)] : $signed(reg54))) && reg17[(1'h1):(1'h0)]) != {$unsigned((reg51[(4'h9):(3'h4)] ?
                      $signed((8'ha7)) : (forvar49 && reg55)))});
            end
          for (forvar57 = (1'h0); (forvar57 < (2'h3)); forvar57 = (forvar57 + (1'h1)))
            begin
              reg58 <= $signed({$signed(($signed(reg43) < (reg55 ?
                      reg23 : forvar47))),
                  (($unsigned(forvar49) == $signed(reg6)) ?
                      {$signed(reg10), $signed(reg55)} : (reg32[(4'hc):(2'h2)] ?
                          reg17 : (^reg54)))});
              reg59 = $unsigned((^reg32));
              reg60 <= $unsigned((forvar47[(2'h3):(2'h3)] - $unsigned((~^forvar47))));
              reg61 <= $unsigned((reg26[(2'h2):(1'h0)] && $unsigned({{forvar57}})));
            end
          reg62 <= reg26[(1'h0):(1'h0)];
        end
    end
  assign wire63 = {$unsigned(reg60), reg55};
  always
    @(posedge clk) begin
      reg64 <= reg45;
      if (reg19)
        begin
          reg65 = reg64;
          reg66 = reg45;
          if ($unsigned($unsigned({$signed((reg37 >>> reg15))})))
            begin
              reg67 = (reg52 ^ ((~$unsigned($signed(reg23))) ?
                  $signed(wire1[(4'h8):(4'h8)]) : reg38));
              reg68 = (~^($signed(reg45[(4'hc):(1'h1)]) ?
                  {{$unsigned((8'hbe))},
                      $signed({reg23})} : reg56[(4'he):(3'h6)]));
              reg69 <= $signed((-{($unsigned(reg15) >>> (reg11 ?
                      reg58 : reg44)),
                  wire0}));
              reg70 <= (reg16 ?
                  (wire2 ?
                      reg61 : (reg52[(4'hb):(1'h0)] >= reg26)) : $unsigned((reg43 * reg26)));
            end
          else
            begin
              reg69 <= ($unsigned(reg66[(1'h0):(1'h0)]) ?
                  $unsigned({(reg26 >>> (wire1 >> wire3))}) : (~|(($unsigned(reg45) ^ (!(8'hb2))) || $unsigned($unsigned((8'hbd))))));
              reg71 = {reg13[(2'h3):(1'h0)],
                  $signed($signed(reg32[(1'h1):(1'h0)]))};
              reg72 <= $unsigned((wire0 + ((~reg29[(2'h2):(1'h0)]) ?
                  (((7'h45) < (8'hbe)) ?
                      (reg44 ? (8'hb8) : wire1) : reg50) : (8'hb9))));
              reg73 = (($signed($signed(((7'h4a) ?
                  reg52 : reg13))) >> ((^~$signed(wire1)) ?
                  (!$unsigned(reg61)) : {wire2,
                      (~^reg10)})) == wire2[(2'h3):(1'h1)]);
              reg74 <= reg17[(3'h4):(2'h3)];
            end
          if ({(~&$signed(reg22))})
            begin
              reg75 <= (^~reg58[(4'h9):(3'h6)]);
              reg76 = ((($unsigned(reg37) ~^ $unsigned((wire4 ?
                          reg50 : reg64))) ?
                      (reg64[(3'h5):(2'h3)] || reg53[(4'he):(3'h4)]) : ($signed($unsigned(reg56)) ?
                          ({reg72, (8'h9c)} ?
                              reg38[(4'hc):(3'h4)] : ((7'h42) ?
                                  reg52 : (8'ha2))) : reg41)) ?
                  $signed($signed((8'hb1))) : (!$signed((wire1 ?
                      $signed(reg61) : $signed(reg55)))));
            end
          else
            begin
              reg75 <= reg72;
              reg77 <= (reg52[(3'h5):(2'h3)] ?
                  $unsigned((~{{reg19}})) : reg16[(2'h3):(2'h3)]);
              reg78 <= ($unsigned((((8'hb2) ^ (reg39 ? reg41 : reg66)) ?
                      reg53 : reg55)) ?
                  (~|(reg39 ~^ ($unsigned(reg60) ?
                      $signed(reg45) : reg38[(3'h4):(1'h0)]))) : $signed($signed(((8'ha4) || reg69[(3'h6):(2'h3)]))));
              reg79 <= reg74[(1'h1):(1'h0)];
              reg80 = $signed(reg15);
            end
        end
      else
        begin
          if ((-reg55))
            begin
              reg69 <= reg72;
            end
          else
            begin
              reg65 = reg11[(2'h3):(1'h1)];
              reg66 = $unsigned((reg77 ?
                  (^~(^$unsigned((8'ha3)))) : (reg78[(4'h9):(1'h0)] ?
                      $signed(reg68) : (((8'hbe) ? reg44 : (8'hba)) ?
                          ((8'h9d) >>> reg30) : reg15))));
              reg67 = wire1;
              reg69 <= reg80[(3'h5):(3'h4)];
            end
          reg70 <= $unsigned(($signed({(reg19 >= reg16), reg71}) ?
              {reg52[(3'h7):(3'h5)],
                  $unsigned(reg71[(4'hb):(4'h8)])} : ($signed($signed(reg55)) ?
                  reg23 : (((8'hb4) ^ reg11) <<< (reg75 ? reg26 : reg23)))));
        end
      for (forvar81 = (1'h0); (forvar81 < (3'h4)); forvar81 = (forvar81 + (1'h1)))
        begin
          reg82 = {(7'h42), reg71[(5'h10):(3'h4)]};
          reg83 = (8'haf);
          for (forvar84 = (1'h0); (forvar84 < (2'h3)); forvar84 = (forvar84 + (1'h1)))
            begin
              reg85 = (((($unsigned(reg19) + reg7) ?
                          reg39 : $unsigned(reg58[(4'h9):(3'h6)])) ?
                      {reg60} : reg41) ?
                  ((^(~|$signed(reg55))) >= reg56) : {$unsigned((+reg82)),
                      {reg74,
                          (((8'hb4) ? reg26 : reg10) ?
                              reg62[(2'h2):(1'h0)] : (reg77 ?
                                  reg19 : reg60))}});
              reg86 = reg32[(1'h0):(1'h0)];
              reg87 <= reg15[(4'h9):(1'h0)];
              reg88 <= $unsigned(($signed(wire2[(2'h2):(1'h1)]) ?
                  $unsigned(((!reg69) && $unsigned(reg32))) : (~|(((8'ha2) ?
                      reg62 : reg43) * (8'ha5)))));
              reg89 <= (~($signed(reg32) >>> wire63));
            end
        end
      if ($signed((^(reg87[(5'h10):(3'h6)] <= (8'h9d)))))
        begin
          for (forvar90 = (1'h0); (forvar90 < (2'h3)); forvar90 = (forvar90 + (1'h1)))
            begin
              reg91 = reg60[(5'h11):(2'h3)];
              reg92 <= (reg80 ?
                  $unsigned((wire4 ?
                      reg61[(4'hf):(1'h0)] : $unsigned(reg60))) : (reg22 ?
                      ({$unsigned(reg53), reg19[(3'h5):(1'h0)]} ?
                          $signed(reg62) : {(~reg87),
                              $unsigned(reg6)}) : (8'hbe)));
              reg93 = (((8'ha2) ?
                      $unsigned($signed((wire0 ?
                          wire2 : reg73))) : $unsigned((-reg64[(4'hd):(3'h4)]))) ?
                  $signed(((^reg74) ?
                      $signed(reg89[(5'h17):(2'h2)]) : (+reg88))) : reg62[(2'h2):(2'h2)]);
              reg94 = $unsigned(reg41);
              reg95 = reg71[(3'h5):(1'h0)];
            end
          reg96 = {(!reg61)};
          reg97 <= reg32;
          if (($unsigned(reg87) * (~^reg69[(1'h0):(1'h0)])))
            begin
              reg98 = {(~^(+$unsigned($unsigned(wire4)))),
                  ((^$unsigned($unsigned(reg43))) < reg16[(2'h2):(2'h2)])};
              reg99 = $signed(reg70[(3'h6):(1'h0)]);
            end
          else
            begin
              reg100 <= (8'hac);
              reg101 = reg80;
              reg102 <= reg15;
              reg103 = $unsigned((|{(8'ha8)}));
              reg104 = $signed(($signed($signed(reg77)) ?
                  (|(~^$signed(reg74))) : $unsigned({(wire63 | reg96),
                      reg96})));
            end
        end
      else
        begin
          reg90 <= (~&$signed(($unsigned($unsigned(reg60)) * reg39[(2'h3):(2'h2)])));
          if ((($signed(reg71) | $signed($signed(reg101[(3'h7):(2'h2)]))) < reg37[(2'h3):(2'h2)]))
            begin
              reg92 <= $signed($signed(reg96[(3'h6):(1'h0)]));
              reg97 <= ($signed((+reg80[(4'ha):(2'h3)])) ?
                  ($unsigned((8'ha3)) ^ $unsigned({(reg97 && reg56),
                      (^~reg62)})) : ((reg73 ?
                      (|(reg80 ?
                          reg97 : (8'ha5))) : (reg37[(3'h6):(3'h4)] << $signed(reg37))) ^ $signed($unsigned({reg19}))));
              reg100 <= reg96[(4'hb):(3'h6)];
              reg101 = $signed(((8'had) + $signed($signed({(8'ha0)}))));
            end
          else
            begin
              reg92 <= $signed((^~{($signed(forvar90) ? (~^reg89) : reg94)}));
              reg97 <= {$signed((|(7'h40)))};
              reg98 = reg100[(2'h2):(2'h2)];
              reg99 = ({reg38[(4'h8):(2'h2)]} ?
                  {($signed($signed(reg79)) ?
                          $unsigned(reg94[(3'h6):(1'h0)]) : $signed((reg41 ~^ reg13)))} : $signed(reg103[(2'h3):(1'h0)]));
              reg100 <= (reg13 ?
                  ((reg60[(5'h12):(3'h5)] ^ $unsigned($signed(reg16))) ?
                      (|(((8'hbe) << reg67) == reg38)) : {(+$signed(reg62))}) : (^wire0[(4'hc):(3'h5)]));
            end
          for (forvar102 = (1'h0); (forvar102 < (2'h3)); forvar102 = (forvar102 + (1'h1)))
            begin
              reg103 = reg44;
            end
          reg105 <= (reg91 ?
              ((^~(~|reg15)) < {((wire2 >>> reg6) ?
                      $unsigned(reg22) : (reg17 ^~ reg50))}) : ({($unsigned(reg50) ?
                      $unsigned(reg72) : (reg83 ? reg100 : reg38)),
                  reg15[(2'h3):(1'h0)]} > (+($signed(reg87) >>> $signed(wire4)))));
          for (forvar106 = (1'h0); (forvar106 < (1'h0)); forvar106 = (forvar106 + (1'h1)))
            begin
              reg107 <= (|{(^reg64)});
              reg108 = reg45;
              reg109 <= $signed(reg74);
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg53)
        begin
          reg110 <= ((reg44[(1'h0):(1'h0)] ?
              (((~^reg60) ? reg30[(5'h16):(4'h9)] : (reg60 ? (7'h4a) : reg87)) ?
                  $signed(reg88[(5'h11):(4'h8)]) : reg61) : $signed(reg19)) >> $signed($signed((8'ha2))));
          reg111 = (|reg30[(4'h8):(2'h3)]);
          for (forvar112 = (1'h0); (forvar112 < (1'h0)); forvar112 = (forvar112 + (1'h1)))
            begin
              reg113 <= reg77[(5'h11):(4'h8)];
              reg114 = ($unsigned($unsigned($signed(((7'h49) + (7'h46))))) ?
                  ($unsigned($signed((~^reg19))) ?
                      wire4[(3'h6):(3'h4)] : wire4) : $signed({reg11}));
              reg115 <= (~&(~(!reg102[(3'h7):(2'h2)])));
              reg116 <= $signed(((~&reg109) ?
                  ((&reg29) ?
                      reg37[(1'h0):(1'h0)] : {reg15,
                          {reg62}}) : (reg113[(4'h8):(3'h7)] ?
                      {reg70[(4'hb):(2'h2)]} : reg97)));
              reg117 <= $unsigned(reg22[(1'h1):(1'h0)]);
            end
          reg118 = reg111;
          if ($unsigned((((!reg37[(3'h6):(3'h6)]) <= $signed({(8'h9c)})) ?
              {(~&$signed(reg62))} : reg38[(1'h1):(1'h1)])))
            begin
              reg119 <= reg117;
              reg120 = {$unsigned(reg97[(4'h9):(2'h2)]), reg17};
              reg121 = (^$unsigned(reg44));
            end
          else
            begin
              reg120 = ($signed(reg26[(1'h1):(1'h0)]) & reg26);
              reg121 = (-wire0[(4'hb):(4'ha)]);
            end
        end
      else
        begin
          reg110 <= reg17;
          for (forvar111 = (1'h0); (forvar111 < (2'h2)); forvar111 = (forvar111 + (1'h1)))
            begin
              reg112 = reg69[(4'hc):(4'hc)];
              reg114 = {reg88,
                  ({{(reg23 ^~ reg114)}, (&$unsigned((7'h44)))} ?
                      (reg114[(1'h1):(1'h0)] ?
                          reg105 : $unsigned((reg11 ?
                              reg43 : wire3))) : ((reg37 < (reg109 && wire63)) ?
                          $signed($unsigned((8'haf))) : reg69))};
              reg115 <= (~^(((7'h43) ?
                  (^~wire63[(2'h2):(2'h2)]) : (^~$unsigned(reg39))) <<< (^({wire1} ?
                  (reg121 ? reg112 : reg50) : $signed((8'hb1))))));
              reg118 = ((&reg26[(2'h2):(2'h2)]) < (8'ha1));
            end
          for (forvar119 = (1'h0); (forvar119 < (2'h3)); forvar119 = (forvar119 + (1'h1)))
            begin
              reg120 = (^($signed((forvar112[(4'hb):(2'h3)] ?
                  $signed(reg113) : (~reg114))) ~^ $signed(($unsigned(reg11) ?
                  (!reg115) : $signed(reg121)))));
            end
          reg122 <= $unsigned(((!reg88) && reg79[(4'hf):(4'hc)]));
          if ((8'h9d))
            begin
              reg123 = (&(reg122 || ({$signed((8'hba))} != ($signed((8'haf)) ?
                  $unsigned(reg110) : (reg113 || (8'hbf))))));
              reg124 = $signed({reg38,
                  (reg111 ?
                      ($signed(reg122) ?
                          reg29 : (reg60 ^~ wire3)) : $signed((!reg53)))});
              reg125 <= (^~$signed(reg38[(3'h7):(3'h5)]));
            end
          else
            begin
              reg125 <= (8'hb9);
              reg126 <= reg45;
              reg127 = (~((8'hae) - reg72[(3'h4):(1'h1)]));
              reg128 = $unsigned((((-$unsigned(reg102)) | (!(-reg61))) ?
                  reg119 : reg30));
            end
        end
      reg129 = $signed(reg109[(2'h2):(2'h2)]);
      if (reg11[(1'h0):(1'h0)])
        begin
          if (((^(!reg79)) > {reg37,
              ({reg39[(1'h1):(1'h0)]} >>> reg114[(1'h1):(1'h0)])}))
            begin
              reg130 <= ($signed({(reg110 >>> ((7'h46) * reg128)),
                  $signed(reg117)}) >= (&reg7[(4'hf):(4'hd)]));
            end
          else
            begin
              reg131 = $unsigned($signed(wire3[(5'h11):(5'h11)]));
              reg132 = ($unsigned($unsigned(reg37[(3'h4):(1'h1)])) ?
                  $unsigned($signed($unsigned(reg114))) : $unsigned((reg16 ?
                      (-$signed(reg88)) : {((8'hb1) ~^ reg7),
                          (reg10 ? reg123 : (8'hb0))})));
              reg133 <= (((reg53 ? reg56 : reg128) ?
                      ($unsigned((~forvar111)) < reg15) : reg44[(4'hd):(2'h2)]) ?
                  $unsigned(reg41) : $signed(reg117[(4'h9):(3'h7)]));
            end
          if (((8'ha2) ?
              (~^$unsigned((~(reg38 << reg132)))) : (~|reg111[(1'h1):(1'h0)])))
            begin
              reg134 <= reg132[(4'hf):(3'h7)];
              reg135 = (&(($signed(reg112) || $unsigned((+(8'ha2)))) ?
                  $signed(reg74) : $unsigned(((reg30 ?
                      (8'hb1) : reg41) && $unsigned((8'ha9))))));
              reg136 <= reg23;
              reg137 = reg50;
              reg138 = reg53;
            end
          else
            begin
              reg135 = $signed(reg38);
              reg136 <= $unsigned(({$signed(((7'h42) ?
                      reg78 : reg29))} >> $unsigned(reg130[(4'he):(4'h8)])));
              reg139 <= wire2;
              reg140 = (~^($signed($signed((-reg138))) + (($unsigned(reg110) || (reg62 || (8'hb7))) ?
                  ($unsigned((8'hbc)) ?
                      ((7'h49) >= (8'ha0)) : $signed(reg111)) : (~^$signed(reg131)))));
            end
          reg141 = {(reg92 | reg130[(3'h5):(2'h2)])};
        end
      else
        begin
          if (reg30[(3'h4):(1'h1)])
            begin
              reg131 = $unsigned((^(^~(|((8'ha9) == wire0)))));
              reg132 = ((!$unsigned(((reg127 & (7'h47)) - ((8'hab) == reg16)))) ?
                  (reg52 ?
                      (|$unsigned($unsigned(reg38))) : reg105) : ((((!reg116) ?
                              (reg90 ? (8'h9c) : reg113) : reg26) ?
                          (|(reg97 ?
                              (8'ha5) : wire4)) : $unsigned($unsigned(reg19))) ?
                      $unsigned(reg127[(1'h0):(1'h0)]) : $signed(reg119)));
              reg133 <= reg77;
            end
          else
            begin
              reg130 <= $unsigned(reg89);
              reg133 <= reg133[(4'h9):(4'h8)];
              reg135 = $unsigned($signed(reg128[(4'hb):(3'h6)]));
            end
        end
      reg142 = $signed($unsigned((~&(+{reg124, reg139}))));
      for (forvar143 = (1'h0); (forvar143 < (1'h1)); forvar143 = (forvar143 + (1'h1)))
        begin
          reg144 = (&{(~|{$signed(reg89), reg17[(4'h9):(3'h4)]}), reg37});
          reg145 <= $signed((^~($signed((reg62 ^ (7'h43))) ?
              ($unsigned(reg124) ? {reg129} : reg26[(2'h2):(1'h1)]) : reg15)));
          for (forvar146 = (1'h0); (forvar146 < (3'h4)); forvar146 = (forvar146 + (1'h1)))
            begin
              reg147 = (~&reg141[(3'h5):(3'h5)]);
              reg148 <= (~&((^(-(reg117 <= reg16))) ~^ reg32[(4'h8):(3'h6)]));
              reg149 = ($signed((|((^~reg117) ?
                  (reg132 << wire3) : $unsigned((8'hbf))))) << $unsigned((|(reg7 ?
                  (reg88 && reg102) : reg130[(4'hf):(1'h1)]))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg150 <= ($unsigned($unsigned(reg107)) * (8'ha3));
      for (forvar151 = (1'h0); (forvar151 < (1'h0)); forvar151 = (forvar151 + (1'h1)))
        begin
          if (reg133)
            begin
              reg152 <= (8'ha1);
              reg153 = $signed($signed(reg117[(4'h8):(3'h7)]));
              reg154 <= reg105[(5'h11):(4'he)];
              reg155 = $signed(reg62[(1'h1):(1'h1)]);
              reg156 <= reg139;
            end
          else
            begin
              reg153 = reg13[(3'h6):(3'h5)];
              reg155 = reg37;
              reg156 <= (+$unsigned($signed(reg58)));
            end
          if (reg115[(3'h5):(1'h1)])
            begin
              reg157 <= reg125;
              reg158 <= $signed((reg97[(4'he):(4'he)] ?
                  {$unsigned(reg152[(2'h2):(1'h1)])} : reg45));
              reg159 <= reg79[(5'h11):(5'h11)];
              reg160 = (8'hb4);
            end
          else
            begin
              reg157 <= (($unsigned({$signed(reg74),
                      $signed(reg125)}) + ((+$unsigned(reg88)) ?
                      ((!reg69) >= {reg56, reg41}) : (!(!reg116)))) ?
                  reg105 : reg72[(4'h9):(1'h1)]);
            end
          reg161 = $signed(reg79);
          reg162 = reg154[(5'h12):(1'h0)];
        end
    end
  always
    @(posedge clk) begin
      reg163 <= $unsigned(((((wire4 ? reg43 : reg44) - reg38[(4'he):(2'h2)]) ?
              (((7'h42) > reg70) - ((8'hae) ?
                  reg7 : reg92)) : ($signed((8'haa)) ? (8'hb3) : reg70)) ?
          ($unsigned(reg45[(4'hd):(4'h9)]) <= reg69) : {$signed(reg159[(3'h4):(2'h2)])}));
    end
  always
    @(posedge clk) begin
      for (forvar164 = (1'h0); (forvar164 < (1'h0)); forvar164 = (forvar164 + (1'h1)))
        begin
          if (($unsigned((reg148 ?
              {reg157[(3'h5):(1'h0)], reg89} : ($signed(reg75) ?
                  $signed(reg39) : reg100[(2'h2):(1'h1)]))) >> (8'h9e)))
            begin
              reg165 <= {reg74, reg22[(1'h1):(1'h1)]};
              reg166 <= reg26;
              reg167 = ($unsigned(reg122) | reg50[(2'h3):(1'h1)]);
              reg168 = reg159;
            end
          else
            begin
              reg167 = reg159[(3'h6):(2'h3)];
            end
          reg169 = $unsigned(reg87[(5'h12):(1'h1)]);
          if ($unsigned({($signed((reg169 << reg52)) ?
                  $signed((reg92 + reg166)) : (((8'h9f) ?
                      reg113 : reg168) > (reg61 ? reg78 : reg58)))}))
            begin
              reg170 <= ($unsigned(reg58) ?
                  $unsigned((+{((7'h41) ? reg50 : reg109)})) : reg38);
              reg171 = ((7'h46) & (wire3 >>> $unsigned(reg148)));
              reg172 <= ((({reg74, (-reg110)} & $signed($signed(reg13))) ?
                      $unsigned(($unsigned((8'h9c)) & (reg92 ?
                          reg58 : reg159))) : ((reg152[(2'h2):(2'h2)] ?
                          (^~reg136) : $signed(reg43)) < $signed((8'ha4)))) ?
                  ($unsigned($unsigned((wire63 ?
                      reg61 : reg29))) <<< ($signed((reg79 != reg150)) ?
                      wire1[(5'h10):(4'hd)] : $signed((~&reg109)))) : reg107);
            end
          else
            begin
              reg170 <= (~&reg52);
              reg171 = ((8'h9c) ?
                  $signed({$unsigned((&wire3))}) : $signed(reg79[(5'h15):(3'h7)]));
              reg172 <= $unsigned(reg72);
            end
          if (((reg77 && $unsigned((~(&reg152)))) ? reg92 : reg75))
            begin
              reg173 = reg158[(3'h5):(1'h0)];
              reg174 = (reg11[(1'h1):(1'h1)] || $signed(reg15));
            end
          else
            begin
              reg173 = reg134;
              reg175 <= ((~(($unsigned(reg17) ~^ reg165) ?
                      (|$unsigned(reg39)) : reg37)) ?
                  reg167[(2'h3):(2'h3)] : (($signed((^~(8'hba))) << reg87) ?
                      ((~{reg60, (8'hbe)}) ?
                          $signed($unsigned((7'h43))) : (^(~&reg60))) : (8'hb7)));
              reg176 = ({wire0[(2'h3):(2'h3)], (7'h43)} ?
                  (((~$unsigned(reg30)) ~^ reg166[(3'h4):(2'h2)]) && ((~^reg45[(3'h5):(2'h2)]) || (reg39 ?
                      (reg130 | reg22) : reg38[(3'h4):(1'h1)]))) : reg15[(2'h3):(2'h3)]);
            end
        end
      reg177 <= {((+$signed($signed(reg22))) ?
              $signed((reg10[(1'h0):(1'h0)] || $unsigned(reg53))) : reg26)};
      for (forvar178 = (1'h0); (forvar178 < (3'h4)); forvar178 = (forvar178 + (1'h1)))
        begin
          reg179 <= (($unsigned(((^reg134) ?
                  (~|reg145) : $signed((8'h9c)))) <= $signed(((forvar164 ?
                      reg109 : wire63) ?
                  $unsigned(reg44) : (8'haa)))) ?
              $unsigned((8'h9f)) : ($signed($signed(reg60[(3'h4):(2'h3)])) ^ (reg39 ?
                  $signed((reg62 ?
                      reg176 : reg117)) : $signed((reg22 - reg150)))));
          reg180 = ((reg41[(1'h0):(1'h0)] ^ $unsigned(reg175)) ?
              (((8'haf) << reg165) ?
                  wire63[(1'h1):(1'h1)] : (reg75 ?
                      reg177[(1'h1):(1'h1)] : $signed((reg176 ?
                          (8'hae) : reg89)))) : $unsigned(((~reg69[(4'hc):(3'h4)]) && (&$unsigned(reg50)))));
          reg181 <= ($signed(reg115) ? reg6 : reg75);
        end
      reg182 <= ($unsigned(reg105[(5'h10):(4'hf)]) && ((reg165 >>> {reg119[(4'hc):(2'h2)]}) > reg64[(4'h8):(3'h6)]));
      reg183 <= (-{$signed(wire3), (^(|$unsigned(wire63)))});
    end
  assign wire184 = $signed((~&({(reg148 ? reg30 : reg10),
                       (|reg77)} <= reg145[(2'h3):(1'h1)])));
  assign wire185 = reg154;
  assign wire186 = reg107[(2'h2):(2'h2)];
  always
    @(posedge clk) begin
      reg187 <= reg157[(3'h6):(2'h3)];
    end
  assign wire188 = (((({reg38} ? $signed((7'h40)) : (!reg64)) ?
                           ({reg122} > ((7'h42) ?
                               reg125 : reg55)) : ($unsigned(reg122) ^ $unsigned(reg16))) ?
                       (8'hbf) : $unsigned(($unsigned(reg105) ?
                           $signed(reg41) : ((7'h47) ?
                               reg19 : reg154)))) == {(8'hac),
                       reg166[(1'h1):(1'h1)]});
  assign wire189 = reg45[(4'h8):(2'h2)];
  assign wire190 = $signed(((reg43 ?
                       (reg107 ?
                           (reg7 ?
                               reg26 : reg105) : (reg79 != reg17)) : ((8'ha9) != $unsigned(reg156))) ^~ ($signed((reg97 ?
                       reg134 : reg148)) <= reg122)));
  always
    @(posedge clk) begin
      reg191 = {reg150};
      if (($unsigned($signed({(reg156 ? reg69 : reg22)})) ?
          reg38[(4'ha):(1'h1)] : reg177[(4'hb):(3'h6)]))
        begin
          reg192 = reg175;
          if ((8'hac))
            begin
              reg193 <= (~|reg23[(3'h4):(1'h1)]);
              reg194 <= {($signed($unsigned($signed(reg55))) ?
                      (8'ha1) : reg115)};
              reg195 <= reg23;
              reg196 <= reg30;
              reg197 <= reg90;
            end
          else
            begin
              reg198 = {(((reg92[(1'h0):(1'h0)] >>> reg197) - $unsigned((-reg44))) >= $unsigned(reg72[(1'h0):(1'h0)])),
                  (7'h45)};
              reg199 <= (reg23[(1'h1):(1'h1)] ?
                  (reg198 ?
                      (reg43 ? reg177 : (^reg38)) : reg16) : {(~&{{reg179},
                          $signed(reg64)})});
            end
          for (forvar200 = (1'h0); (forvar200 < (1'h1)); forvar200 = (forvar200 + (1'h1)))
            begin
              reg201 <= (8'ha4);
              reg202 <= reg56;
              reg203 <= {reg97, reg148};
              reg204 = $unsigned($unsigned(((reg198[(1'h1):(1'h0)] ^ (reg156 >> reg136)) ?
                  (reg109 - (+reg88)) : $signed((reg45 ? reg69 : reg26)))));
              reg205 <= $signed((^~{($unsigned(reg10) > wire184[(4'hd):(4'h8)])}));
            end
        end
      else
        begin
          reg193 <= reg159[(4'hf):(4'hf)];
          for (forvar194 = (1'h0); (forvar194 < (2'h2)); forvar194 = (forvar194 + (1'h1)))
            begin
              reg198 = (&reg38);
              reg199 <= reg203;
              reg200 = $unsigned((+(8'ha7)));
              reg204 = {{(!$unsigned((reg55 + (7'h40))))},
                  $signed(wire4[(2'h3):(1'h1)])};
              reg205 <= (~|{($unsigned((reg58 == reg200)) ?
                      reg115 : (^(reg43 * reg199))),
                  $signed(reg198)});
            end
          reg206 <= (-(8'hae));
          for (forvar207 = (1'h0); (forvar207 < (1'h0)); forvar207 = (forvar207 + (1'h1)))
            begin
              reg208 <= (((~|$signed(reg100[(2'h3):(1'h0)])) <<< reg165) <<< $signed((reg56 || ((reg15 ?
                  (7'h47) : reg159) == reg191))));
              reg209 = (8'ha2);
              reg210 = (~({$unsigned((forvar200 != reg64)), (|(^~reg126))} ?
                  ($signed((reg126 ?
                      reg64 : reg125)) + $signed((8'ha8))) : ($unsigned($signed(wire188)) || reg6[(1'h0):(1'h0)])));
            end
        end
      reg211 = reg203;
      reg212 <= reg163;
      for (forvar213 = (1'h0); (forvar213 < (2'h2)); forvar213 = (forvar213 + (1'h1)))
        begin
          reg214 <= reg159[(5'h11):(4'he)];
          reg215 <= ((^~reg133) ?
              $unsigned((reg214[(1'h1):(1'h0)] >> $unsigned(reg195[(2'h2):(1'h0)]))) : (reg69 | reg75[(1'h1):(1'h1)]));
          for (forvar216 = (1'h0); (forvar216 < (2'h2)); forvar216 = (forvar216 + (1'h1)))
            begin
              reg217 <= $signed(reg194[(3'h4):(1'h0)]);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar218 = (1'h0); (forvar218 < (3'h4)); forvar218 = (forvar218 + (1'h1)))
        begin
          reg219 = (+({($signed(reg19) ^~ $signed(reg195)),
              $signed((-reg197))} >= (reg74[(3'h6):(3'h4)] ?
              $unsigned({(7'h40)}) : (-(8'h9c)))));
          reg220 <= $signed(($unsigned((reg88 ?
              $unsigned((8'hac)) : reg165)) << reg116));
          for (forvar221 = (1'h0); (forvar221 < (2'h2)); forvar221 = (forvar221 + (1'h1)))
            begin
              reg222 = wire0;
              reg223 <= reg50[(4'ha):(4'ha)];
              reg224 = reg177;
              reg225 = ($unsigned($signed(reg19)) ?
                  ((^$unsigned(reg44[(4'hc):(4'h9)])) == $unsigned(reg158)) : reg133[(3'h7):(2'h2)]);
              reg226 = ((~|$unsigned(reg195[(4'h8):(3'h7)])) ?
                  (~^$unsigned(reg105[(4'h9):(3'h5)])) : $unsigned($unsigned(reg74)));
            end
          for (forvar227 = (1'h0); (forvar227 < (2'h2)); forvar227 = (forvar227 + (1'h1)))
            begin
              reg228 <= (~&reg179);
              reg229 <= reg166;
              reg230 = $unsigned($unsigned($signed($unsigned(wire190[(2'h2):(1'h1)]))));
              reg231 <= reg203[(4'he):(4'hd)];
            end
          for (forvar232 = (1'h0); (forvar232 < (1'h1)); forvar232 = (forvar232 + (1'h1)))
            begin
              reg233 = reg228;
              reg234 = reg100;
              reg235 <= reg88;
              reg236 = $unsigned($unsigned($unsigned(($unsigned(forvar218) ?
                  (^~reg122) : (~^forvar221)))));
            end
        end
      for (forvar237 = (1'h0); (forvar237 < (3'h4)); forvar237 = (forvar237 + (1'h1)))
        begin
          reg238 = reg228;
          for (forvar239 = (1'h0); (forvar239 < (1'h1)); forvar239 = (forvar239 + (1'h1)))
            begin
              reg240 <= $signed(forvar221);
              reg241 <= (($unsigned($signed($unsigned(reg166))) >= $unsigned((+$unsigned(reg223)))) ?
                  ((~^$unsigned((~reg44))) ?
                      $signed(reg102) : (~^wire63)) : $unsigned(reg215[(2'h2):(1'h0)]));
              reg242 = wire3;
              reg243 = (+reg226[(2'h3):(1'h0)]);
              reg244 = ({(+$signed((reg6 ? reg238 : wire4))),
                  $signed((~$signed((7'h47))))} - (~((~^$signed(reg29)) ?
                  $signed(reg154[(4'h8):(4'h8)]) : (~{reg75, reg52}))));
            end
          if ($unsigned(reg224))
            begin
              reg245 = ($signed($signed(((forvar218 ?
                  (8'hbf) : wire4) | (~&reg41)))) != (reg238 ?
                  (reg226 | (7'h41)) : $unsigned(reg136[(5'h17):(4'hb)])));
              reg246 <= ($unsigned($unsigned($unsigned((~|reg7)))) ?
                  $unsigned(reg199[(3'h7):(3'h5)]) : $unsigned({forvar237[(1'h0):(1'h0)],
                      ($unsigned(wire185) ?
                          reg32[(4'h8):(4'h8)] : $signed((8'ha8)))}));
              reg247 <= ((^(~^(&(reg215 ^~ reg224)))) >= ($unsigned((reg23 ?
                      reg217 : reg243[(2'h3):(2'h2)])) ?
                  ((-$signed(forvar239)) ?
                      reg182 : ((reg165 & reg202) <<< (&(7'h48)))) : $unsigned(($unsigned(reg197) ?
                      reg69 : $signed(wire1)))));
              reg248 <= (~^reg22);
            end
          else
            begin
              reg246 <= $signed(wire185[(4'he):(2'h3)]);
              reg247 <= (~|($unsigned(reg37[(3'h6):(1'h1)]) || $unsigned($signed($unsigned(reg69)))));
              reg249 = $unsigned($signed($unsigned({reg130[(4'hc):(1'h0)]})));
              reg250 = ($signed(reg172[(3'h6):(3'h5)]) ?
                  {reg150[(2'h2):(1'h0)]} : reg16);
              reg251 = $signed($unsigned(((-reg222) ^ reg53)));
            end
          reg252 = ($signed($signed((^(~^(8'ha5))))) >= $unsigned(((reg115[(4'h9):(2'h2)] ?
                  $signed(reg215) : (8'h9f)) ?
              (^$unsigned((8'had))) : ((reg163 + reg29) >>> reg187))));
          if (reg240)
            begin
              reg253 = (({reg126[(2'h3):(2'h3)]} > $unsigned(((reg157 * reg224) && (reg116 ?
                  reg126 : reg166)))) & {$unsigned(((reg126 ?
                      reg235 : reg220) <= $unsigned(reg163))),
                  $signed({(^~reg41)})});
              reg254 = ($unsigned((($signed(reg226) <= reg16) & $signed((forvar237 ?
                      reg43 : reg238)))) ?
                  $unsigned(($unsigned(forvar237[(1'h1):(1'h1)]) < ($signed((8'hbe)) ?
                      $unsigned(reg154) : {reg75}))) : (!($signed((reg148 > reg75)) ?
                      reg219 : $signed({reg248}))));
              reg255 <= (-reg226[(2'h2):(1'h1)]);
            end
          else
            begin
              reg253 = $unsigned((((~(reg212 ?
                      reg13 : reg226)) & $unsigned((reg208 != reg172))) ?
                  {{$unsigned(wire2), reg194}} : $signed(reg215)));
              reg254 = (~&(8'hb1));
              reg256 = ((reg195 ?
                  $signed((reg70[(4'h8):(3'h6)] ?
                      (~&reg215) : (reg102 <= reg107))) : (~&reg79)) << (reg10[(1'h0):(1'h0)] ?
                  $signed(((reg115 ?
                      reg6 : reg38) < reg53[(4'hc):(3'h4)])) : $unsigned((^{reg255}))));
            end
        end
      if ((^(($unsigned((reg251 ? reg64 : reg244)) ?
          ($signed(reg154) > (&reg38)) : $signed((reg89 ?
              wire186 : reg205))) - reg249)))
        begin
          if ($signed((8'haa)))
            begin
              reg257 = $signed(wire0[(3'h4):(1'h1)]);
              reg258 <= $unsigned((~{((-reg248) >> (reg187 - reg166))}));
              reg259 = $unsigned((+(reg61 ?
                  ($unsigned((8'hb4)) == (~^(8'hac))) : ((reg170 == reg62) ?
                      ((7'h47) <<< reg159) : reg199[(2'h3):(2'h2)]))));
              reg260 <= reg156;
              reg261 = reg229;
            end
          else
            begin
              reg257 = reg247;
            end
          reg262 <= (((((reg56 != reg130) <<< (8'hbd)) | (reg236 ^~ reg56[(4'hc):(4'ha)])) | wire186) >>> $signed((-reg158)));
        end
      else
        begin
          for (forvar257 = (1'h0); (forvar257 < (2'h2)); forvar257 = (forvar257 + (1'h1)))
            begin
              reg258 <= ((-reg172) != {$signed($unsigned($signed(forvar232)))});
              reg259 = $signed((($unsigned((reg97 >> (8'h9f))) ?
                      (|reg126) : reg150) ?
                  (((reg29 ? reg37 : reg187) ?
                          $signed(reg32) : $signed(reg175)) ?
                      ($signed(reg70) ?
                          (7'h49) : (reg219 <= reg202)) : ((^~reg205) ?
                          (wire190 ?
                              reg102 : reg245) : $signed(reg105))) : ((~(&reg117)) == $unsigned(((8'hb6) < reg228)))));
            end
          reg261 = {(reg150 ?
                  $signed(reg22[(2'h2):(1'h1)]) : (((|reg58) ?
                      reg233[(3'h5):(2'h2)] : reg157[(3'h4):(2'h2)]) - (forvar257[(4'h8):(1'h1)] != {wire4,
                      reg195})))};
          reg263 = $unsigned($unsigned($unsigned(reg252)));
          for (forvar264 = (1'h0); (forvar264 < (2'h2)); forvar264 = (forvar264 + (1'h1)))
            begin
              reg265 = ($unsigned((|$signed(((8'h9e) ^~ reg197)))) <= reg199);
              reg266 = (reg154 ?
                  (~&reg90[(1'h1):(1'h1)]) : ($signed((reg254[(4'hf):(4'hc)] ?
                      $signed(reg238) : (reg236 ?
                          forvar232 : (8'ha0)))) - {((reg16 >>> reg77) ?
                          (reg217 ~^ reg119) : wire4[(3'h5):(3'h4)])}));
            end
          for (forvar267 = (1'h0); (forvar267 < (1'h1)); forvar267 = (forvar267 + (1'h1)))
            begin
              reg268 <= (($unsigned(((+reg220) > (reg197 ? reg222 : reg89))) ?
                  $signed({$signed(reg233)}) : $unsigned((~&(~|reg195)))) - $signed($unsigned($unsigned((^reg222)))));
              reg269 = $unsigned($signed($signed($signed($unsigned((7'h49))))));
            end
        end
    end
  assign wire270 = ($signed($unsigned($signed((reg187 && reg150)))) ?
                       $signed((~|reg205)) : (reg165[(5'h11):(1'h0)] | $unsigned(((reg64 ?
                               reg154 : reg87) ?
                           $unsigned(reg90) : (|reg37)))));
  assign wire271 = reg50[(3'h7):(2'h3)];
  assign wire272 = (((^~((reg223 <= reg220) ?
                           (reg102 << reg136) : $unsigned((7'h42)))) - $unsigned($signed({wire188,
                           reg170}))) ?
                       (wire184[(5'h12):(4'hf)] << $unsigned($signed(wire63[(4'h9):(4'h8)]))) : (~|((~^{reg58}) ?
                           (reg199 ?
                               wire0[(3'h5):(3'h4)] : reg133[(3'h6):(3'h6)]) : reg62)));
  module273 #() modinst1468 (wire1467, clk, reg215, reg50, reg165, wire2, wire4);
  always
    @(posedge clk) begin
      reg1469 = reg203[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg1470 = (($unsigned(reg58[(1'h0):(1'h0)]) >> $unsigned(((reg260 >> reg44) << $signed(reg262)))) <<< (~$signed((reg181 ?
          $unsigned(reg154) : (reg41 ? wire270 : reg60)))));
      if ($signed(reg208))
        begin
          if ($unsigned(((({reg102, (8'haf)} * (reg89 ^~ reg109)) ?
                  $unsigned($signed(reg107)) : (~^$unsigned(wire270))) ?
              $unsigned({(reg79 - reg107)}) : (reg116[(3'h5):(1'h0)] <= $unsigned({wire270})))))
            begin
              reg1471 <= $signed((8'had));
              reg1472 <= reg43;
              reg1473 <= (+{reg152[(1'h1):(1'h1)]});
            end
          else
            begin
              reg1474 = $unsigned($signed((7'h45)));
              reg1475 <= (~&(~$unsigned(({reg109} <= $signed(reg170)))));
              reg1476 = (~^{(~|$unsigned($unsigned(wire63))),
                  {reg182, $unsigned(reg187)}});
              reg1477 = $signed($signed((reg1473 ?
                  {wire272[(4'h9):(3'h5)], (reg248 * reg181)} : reg60)));
            end
          reg1478 = $unsigned($unsigned($signed($unsigned((-reg6)))));
          reg1479 <= $signed(reg52);
          if ((reg62[(1'h1):(1'h1)] ?
              reg268 : (((reg170[(5'h17):(3'h6)] ?
                          reg260[(4'hb):(4'ha)] : (reg89 ? reg255 : reg1477)) ?
                      ($signed(wire186) <= (reg13 >> reg92)) : ((reg208 ?
                              reg87 : (8'hbd)) ?
                          (+reg165) : {reg19, reg64})) ?
                  ((~reg196[(2'h3):(2'h3)]) ?
                      reg45 : $signed($unsigned((7'h40)))) : $signed($unsigned(reg159)))))
            begin
              reg1480 <= reg16[(3'h6):(1'h0)];
              reg1481 <= (~|{$signed({((8'ha0) ? wire272 : reg202), (7'h47)})});
              reg1482 = reg88;
              reg1483 = {((^(^~reg52)) ?
                      $signed(reg175) : reg154[(3'h4):(1'h1)])};
            end
          else
            begin
              reg1482 = reg11;
              reg1484 <= (reg58 ? reg220 : reg268);
              reg1485 <= $unsigned($unsigned(($signed($signed(reg228)) && reg247)));
              reg1486 = reg10[(3'h7):(1'h0)];
            end
        end
      else
        begin
          if (((($signed((~^(8'hb5))) ?
              ($signed(wire272) ?
                  (wire3 && reg177) : reg1483) : $signed($unsigned(reg89))) <<< $unsigned(((reg92 ?
                  reg1486 : (8'ha5)) ?
              $signed(reg134) : ((8'hb7) ?
                  reg1474 : reg199)))) >>> $unsigned($unsigned((~|reg1484)))))
            begin
              reg1474 = $signed((&reg1481[(4'hd):(2'h2)]));
              reg1476 = (+($signed($signed(((8'hb5) ?
                  reg22 : reg6))) + (reg50 >= $unsigned($signed(reg157)))));
              reg1477 = (reg235[(1'h0):(1'h0)] ~^ (+reg170[(4'h9):(2'h2)]));
              reg1479 <= $signed(reg181);
              reg1482 = ((reg214[(1'h0):(1'h0)] ?
                      $unsigned($signed((~&wire0))) : $unsigned(reg148)) ?
                  (($unsigned($signed(reg26)) ^ reg229[(4'ha):(4'h9)]) ^ reg262[(4'ha):(2'h2)]) : reg105);
            end
          else
            begin
              reg1471 <= (|(~((|reg159) >= $unsigned(reg45))));
              reg1472 <= ((((reg159 ? {reg1476, reg15} : (^~reg1471)) ?
                      $signed((reg38 & reg217)) : {wire188}) != ($unsigned($unsigned(wire0)) > ({reg255} ?
                      (8'hb3) : (reg72 ? reg177 : reg1481)))) ?
                  (reg240[(1'h0):(1'h0)] ?
                      reg53[(4'he):(4'hb)] : (reg228 ~^ ((reg29 <<< reg1472) && (reg38 ~^ reg196)))) : reg163[(1'h0):(1'h0)]);
              reg1473 <= (reg156 << (7'h4a));
              reg1474 = reg11[(2'h2):(2'h2)];
            end
          reg1483 = reg16[(3'h6):(3'h6)];
          if (reg50)
            begin
              reg1486 = $unsigned({$unsigned($signed((8'ha8)))});
              reg1487 <= $signed((|($unsigned({reg1480}) ?
                  $signed(reg193[(1'h0):(1'h0)]) : reg1476)));
              reg1488 <= $unsigned($signed((((~|reg39) ^ (reg29 ?
                      reg1477 : (7'h40))) ?
                  (reg229 ?
                      (~^(8'hbf)) : reg56[(5'h10):(4'hb)]) : $signed($signed(reg156)))));
            end
          else
            begin
              reg1486 = reg17[(1'h0):(1'h0)];
            end
          reg1489 <= ((~|(8'ha3)) ? (7'h41) : reg154[(4'hf):(3'h5)]);
          if ((($signed(($signed(reg1481) >>> $unsigned(reg255))) ?
              (|{(reg182 ? reg16 : reg44),
                  (reg69 | wire4)}) : ((^(reg182 & (8'hb1))) ?
                  $signed(reg44[(4'he):(4'hd)]) : (((8'ha4) >> reg134) > $signed((8'ha4))))) << reg170))
            begin
              reg1490 = (((+{reg39, (reg248 ? reg159 : (7'h4a))}) ?
                  $unsigned(((reg1487 == reg102) ?
                      (wire1 ?
                          (8'hba) : (7'h46)) : (~|reg196))) : ($signed(reg1484) && (~^reg113[(3'h7):(1'h1)]))) - {{reg89[(4'hc):(4'hc)]}});
              reg1491 = reg134;
            end
          else
            begin
              reg1490 = $signed((wire272 - reg29[(1'h0):(1'h0)]));
              reg1491 = reg1491;
            end
        end
    end
  assign wire1492 = $unsigned({reg70, (~&(~(wire186 ? reg240 : reg16)))});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module273  (y, clk, wire274, wire275, wire276, wire277, wire278);
  output wire [(32'hb2d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h16):(1'h0)] wire274;
  input wire signed [(5'h11):(1'h0)] wire275;
  input wire signed [(4'he):(1'h0)] wire276;
  input wire [(5'h15):(1'h0)] wire277;
  input wire signed [(5'h11):(1'h0)] wire278;
  wire signed [(4'he):(1'h0)] wire1453;
  wire [(3'h6):(1'h0)] wire1411;
  wire [(5'h14):(1'h0)] wire1315;
  wire [(5'h17):(1'h0)] wire668;
  wire signed [(5'h10):(1'h0)] wire653;
  wire [(4'hb):(1'h0)] wire652;
  wire [(5'h18):(1'h0)] wire650;
  wire signed [(5'h16):(1'h0)] wire1317;
  wire [(2'h2):(1'h0)] wire1345;
  wire signed [(4'h8):(1'h0)] wire1346;
  wire [(5'h10):(1'h0)] wire1409;
  reg [(4'hb):(1'h0)] reg1464 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1463 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1461 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1460 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1458 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1457 = (1'h0);
  reg [(4'hc):(1'h0)] reg1455 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1408 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1407 = (1'h0);
  reg [(4'hd):(1'h0)] reg1405 = (1'h0);
  reg [(5'h11):(1'h0)] reg1404 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1399 = (1'h0);
  reg [(5'h11):(1'h0)] reg1396 = (1'h0);
  reg [(4'hf):(1'h0)] reg1395 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1393 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1387 = (1'h0);
  reg [(3'h4):(1'h0)] reg1386 = (1'h0);
  reg [(4'ha):(1'h0)] reg1383 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1381 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1378 = (1'h0);
  reg [(5'h16):(1'h0)] reg1377 = (1'h0);
  reg [(5'h16):(1'h0)] reg1374 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1373 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1372 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1370 = (1'h0);
  reg [(3'h6):(1'h0)] reg1369 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1367 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1366 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1365 = (1'h0);
  reg [(5'h15):(1'h0)] reg1363 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1360 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1357 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1355 = (1'h0);
  reg [(5'h12):(1'h0)] reg1352 = (1'h0);
  reg [(3'h4):(1'h0)] reg1350 = (1'h0);
  reg [(2'h3):(1'h0)] reg1349 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1348 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1347 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1343 = (1'h0);
  reg [(3'h7):(1'h0)] reg1342 = (1'h0);
  reg [(5'h13):(1'h0)] reg1340 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1339 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1338 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1335 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1334 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1333 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1331 = (1'h0);
  reg [(5'h16):(1'h0)] reg1330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1329 = (1'h0);
  reg [(5'h15):(1'h0)] reg1327 = (1'h0);
  reg [(5'h16):(1'h0)] reg1325 = (1'h0);
  reg [(5'h17):(1'h0)] reg1323 = (1'h0);
  reg [(4'h8):(1'h0)] reg1319 = (1'h0);
  reg [(5'h16):(1'h0)] reg658 = (1'h0);
  reg [(3'h6):(1'h0)] reg661 = (1'h0);
  reg [(3'h5):(1'h0)] reg663 = (1'h0);
  reg [(4'ha):(1'h0)] reg666 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg667 = (1'h0);
  reg [(5'h11):(1'h0)] reg670 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg671 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg674 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg675 = (1'h0);
  reg [(5'h18):(1'h0)] reg676 = (1'h0);
  reg [(5'h16):(1'h0)] reg678 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg679 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg683 = (1'h0);
  reg [(5'h10):(1'h0)] reg684 = (1'h0);
  reg [(5'h14):(1'h0)] reg685 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg691 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg692 = (1'h0);
  reg signed [(4'he):(1'h0)] reg693 = (1'h0);
  reg [(4'hf):(1'h0)] reg695 = (1'h0);
  reg [(3'h6):(1'h0)] reg697 = (1'h0);
  reg signed [(4'he):(1'h0)] reg699 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg702 = (1'h0);
  reg [(5'h13):(1'h0)] reg1415 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1416 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1417 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1420 = (1'h0);
  reg [(5'h15):(1'h0)] reg1421 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1422 = (1'h0);
  reg [(4'hd):(1'h0)] reg1423 = (1'h0);
  reg [(4'hf):(1'h0)] reg1424 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1428 = (1'h0);
  reg [(4'h8):(1'h0)] reg1431 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1433 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1434 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1435 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1437 = (1'h0);
  reg [(5'h16):(1'h0)] reg1438 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1442 = (1'h0);
  reg [(2'h3):(1'h0)] reg1444 = (1'h0);
  reg [(4'he):(1'h0)] reg1446 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1449 = (1'h0);
  reg [(5'h10):(1'h0)] reg1451 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1466 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1465 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1462 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1459 = (1'h0);
  reg [(5'h16):(1'h0)] forvar1456 = (1'h0);
  reg [(5'h13):(1'h0)] reg1452 = (1'h0);
  reg [(5'h12):(1'h0)] reg1450 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1448 = (1'h0);
  reg [(5'h10):(1'h0)] reg1447 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1445 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1443 = (1'h0);
  reg [(5'h10):(1'h0)] reg1441 = (1'h0);
  reg [(4'hb):(1'h0)] reg1440 = (1'h0);
  reg [(4'ha):(1'h0)] reg1439 = (1'h0);
  reg [(5'h18):(1'h0)] reg1436 = (1'h0);
  reg [(4'he):(1'h0)] reg1432 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1430 = (1'h0);
  reg [(4'hb):(1'h0)] reg1429 = (1'h0);
  reg [(5'h10):(1'h0)] reg1427 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1426 = (1'h0);
  reg [(5'h14):(1'h0)] reg1425 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1419 = (1'h0);
  reg [(5'h15):(1'h0)] reg1418 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1414 = (1'h0);
  reg [(4'hb):(1'h0)] reg1413 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1406 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1403 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1402 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1401 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1400 = (1'h0);
  reg [(4'hd):(1'h0)] reg1398 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1397 = (1'h0);
  reg [(3'h7):(1'h0)] reg1394 = (1'h0);
  reg [(5'h13):(1'h0)] reg1392 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1391 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1390 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1389 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1388 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1385 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1384 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1382 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1380 = (1'h0);
  reg [(5'h17):(1'h0)] reg1379 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1378 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1376 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1375 = (1'h0);
  reg [(4'hf):(1'h0)] reg1371 = (1'h0);
  reg [(3'h4):(1'h0)] reg1368 = (1'h0);
  reg [(4'hb):(1'h0)] reg1364 = (1'h0);
  reg [(4'he):(1'h0)] forvar1362 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1361 = (1'h0);
  reg [(3'h7):(1'h0)] reg1359 = (1'h0);
  reg [(4'hf):(1'h0)] reg1358 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar1353 = (1'h0);
  reg [(4'ha):(1'h0)] reg1356 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1354 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1353 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1351 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1344 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar1341 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1337 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1336 = (1'h0);
  reg [(5'h15):(1'h0)] reg1332 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1328 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1326 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1324 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1322 = (1'h0);
  reg [(4'hc):(1'h0)] reg1321 = (1'h0);
  reg [(4'h8):(1'h0)] reg1320 = (1'h0);
  reg [(2'h2):(1'h0)] reg701 = (1'h0);
  reg signed [(4'he):(1'h0)] reg700 = (1'h0);
  reg [(3'h7):(1'h0)] reg698 = (1'h0);
  reg [(5'h12):(1'h0)] reg696 = (1'h0);
  reg [(2'h3):(1'h0)] reg694 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg690 = (1'h0);
  reg [(4'hc):(1'h0)] reg689 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar688 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg687 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg686 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar682 = (1'h0);
  reg [(2'h2):(1'h0)] reg681 = (1'h0);
  reg [(3'h7):(1'h0)] reg680 = (1'h0);
  reg [(5'h12):(1'h0)] reg677 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg673 = (1'h0);
  reg [(4'hb):(1'h0)] reg672 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar669 = (1'h0);
  reg [(5'h16):(1'h0)] reg662 = (1'h0);
  reg [(4'h8):(1'h0)] reg665 = (1'h0);
  reg [(4'hf):(1'h0)] reg664 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar662 = (1'h0);
  reg [(5'h12):(1'h0)] reg660 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar659 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg657 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg656 = (1'h0);
  reg [(3'h4):(1'h0)] reg655 = (1'h0);
  reg [(2'h2):(1'h0)] forvar654 = (1'h0);
  assign y = {wire1453,
                 wire1411,
                 wire1315,
                 wire668,
                 wire653,
                 wire652,
                 wire650,
                 wire1317,
                 wire1345,
                 wire1346,
                 wire1409,
                 reg1464,
                 reg1463,
                 reg1461,
                 reg1460,
                 reg1458,
                 reg1457,
                 reg1455,
                 reg1408,
                 reg1407,
                 reg1405,
                 reg1404,
                 reg1399,
                 reg1396,
                 reg1395,
                 reg1393,
                 reg1387,
                 reg1386,
                 reg1383,
                 reg1381,
                 reg1378,
                 reg1377,
                 reg1374,
                 reg1373,
                 reg1372,
                 reg1370,
                 reg1369,
                 reg1367,
                 reg1366,
                 reg1365,
                 reg1363,
                 reg1360,
                 reg1357,
                 reg1355,
                 reg1352,
                 reg1350,
                 reg1349,
                 reg1348,
                 reg1347,
                 reg1343,
                 reg1342,
                 reg1340,
                 reg1339,
                 reg1338,
                 reg1335,
                 reg1334,
                 reg1333,
                 reg1331,
                 reg1330,
                 reg1329,
                 reg1327,
                 reg1325,
                 reg1323,
                 reg1319,
                 reg658,
                 reg661,
                 reg663,
                 reg666,
                 reg667,
                 reg670,
                 reg671,
                 reg674,
                 reg675,
                 reg676,
                 reg678,
                 reg679,
                 reg683,
                 reg684,
                 reg685,
                 reg691,
                 reg692,
                 reg693,
                 reg695,
                 reg697,
                 reg699,
                 reg702,
                 reg1415,
                 reg1416,
                 reg1417,
                 reg1420,
                 reg1421,
                 reg1422,
                 reg1423,
                 reg1424,
                 reg1428,
                 reg1431,
                 reg1433,
                 reg1434,
                 reg1435,
                 reg1437,
                 reg1438,
                 reg1442,
                 reg1444,
                 reg1446,
                 reg1449,
                 reg1451,
                 reg1466,
                 reg1465,
                 forvar1462,
                 reg1459,
                 forvar1456,
                 reg1452,
                 reg1450,
                 forvar1448,
                 reg1447,
                 forvar1445,
                 forvar1443,
                 reg1441,
                 reg1440,
                 reg1439,
                 reg1436,
                 reg1432,
                 forvar1430,
                 reg1429,
                 reg1427,
                 reg1426,
                 reg1425,
                 reg1419,
                 reg1418,
                 forvar1414,
                 reg1413,
                 reg1406,
                 forvar1403,
                 forvar1402,
                 reg1401,
                 forvar1400,
                 reg1398,
                 reg1397,
                 reg1394,
                 reg1392,
                 reg1391,
                 reg1390,
                 reg1389,
                 forvar1388,
                 forvar1385,
                 reg1384,
                 reg1382,
                 reg1380,
                 reg1379,
                 forvar1378,
                 reg1376,
                 reg1375,
                 reg1371,
                 reg1368,
                 reg1364,
                 forvar1362,
                 forvar1361,
                 reg1359,
                 reg1358,
                 forvar1353,
                 reg1356,
                 reg1354,
                 reg1353,
                 reg1351,
                 reg1344,
                 forvar1341,
                 forvar1337,
                 reg1336,
                 reg1332,
                 reg1328,
                 reg1326,
                 forvar1324,
                 forvar1322,
                 reg1321,
                 reg1320,
                 reg701,
                 reg700,
                 reg698,
                 reg696,
                 reg694,
                 reg690,
                 reg689,
                 forvar688,
                 reg687,
                 reg686,
                 forvar682,
                 reg681,
                 reg680,
                 reg677,
                 reg673,
                 reg672,
                 forvar669,
                 reg662,
                 reg665,
                 reg664,
                 forvar662,
                 reg660,
                 forvar659,
                 reg657,
                 reg656,
                 reg655,
                 forvar654,
                 (1'h0)};
  module279 #() modinst651 (.wire281(wire277), .wire280(wire278), .y(wire650), .wire284(wire275), .wire282(wire276), .clk(clk), .wire283(wire274));
  assign wire652 = wire275;
  assign wire653 = ((|{((wire650 ? wire276 : wire650) ?
                               ((8'hba) ?
                                   wire274 : (8'hbf)) : (wire652 >>> wire274)),
                           wire276[(3'h4):(2'h2)]}) ?
                       (+(&(wire652 ~^ (wire278 == wire650)))) : $signed((wire652[(3'h6):(2'h2)] ?
                           ((wire276 + wire650) || (+wire278)) : $unsigned(wire652))));
  always
    @(posedge clk) begin
      for (forvar654 = (1'h0); (forvar654 < (2'h2)); forvar654 = (forvar654 + (1'h1)))
        begin
          reg655 = {(wire652 ^~ wire275[(4'hd):(1'h0)])};
        end
      reg656 = wire274;
      reg657 = {($unsigned(reg656[(4'hf):(3'h6)]) && (forvar654[(2'h2):(1'h0)] ?
              wire278 : $unsigned($signed(reg655)))),
          (^~wire274)};
      reg658 <= $signed(({wire278[(4'hd):(4'hb)],
              ((^~forvar654) << {(8'ha4), wire275})} ?
          wire652[(2'h2):(1'h0)] : (&$signed(((8'haa) | reg655)))));
    end
  always
    @(posedge clk) begin
      if ($signed(wire277))
        begin
          for (forvar659 = (1'h0); (forvar659 < (1'h1)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 = $signed($unsigned($unsigned(wire650[(4'hf):(4'hc)])));
            end
          reg661 <= (^~wire276[(4'he):(4'h9)]);
          for (forvar662 = (1'h0); (forvar662 < (2'h2)); forvar662 = (forvar662 + (1'h1)))
            begin
              reg663 <= reg661[(2'h3):(2'h3)];
              reg664 = reg661[(2'h3):(2'h3)];
              reg665 = $unsigned(((&reg664) != $signed($unsigned((-(8'hbc))))));
            end
        end
      else
        begin
          for (forvar659 = (1'h0); (forvar659 < (2'h3)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 = $signed($unsigned(($unsigned((|wire653)) ?
                  reg661 : $unsigned((reg663 ? wire650 : wire653)))));
              reg662 = (~|forvar662[(1'h0):(1'h0)]);
            end
          reg664 = reg660;
          reg665 = $unsigned({(wire277 ^ {$signed((8'hb6))})});
        end
      reg666 <= reg664;
      reg667 <= (^~((($unsigned(wire653) - $signed(forvar662)) ?
          ((wire275 ? reg666 : forvar662) ?
              {reg666} : $signed(wire276)) : (&forvar662[(5'h14):(3'h4)])) && (($unsigned(forvar659) ?
              {reg661} : (reg666 ? reg660 : reg665)) ?
          wire278 : ((wire650 ? forvar659 : forvar659) ?
              (reg661 ? (8'ha2) : (8'hab)) : reg666[(1'h1):(1'h0)]))));
    end
  assign wire668 = (+(-wire650[(3'h6):(3'h6)]));
  always
    @(posedge clk) begin
      for (forvar669 = (1'h0); (forvar669 < (1'h0)); forvar669 = (forvar669 + (1'h1)))
        begin
          reg670 <= (reg658[(3'h7):(3'h7)] >= $signed(wire650));
          if ($signed(wire278))
            begin
              reg671 <= $unsigned((~(~wire652[(3'h5):(1'h0)])));
              reg672 = wire668[(1'h1):(1'h1)];
              reg673 = (!wire652);
            end
          else
            begin
              reg672 = (((reg663 ?
                      ($unsigned(forvar669) ?
                          (reg672 ~^ reg663) : $signed(reg663)) : (+$unsigned(wire278))) != ($signed($signed(reg666)) ?
                      (8'hbd) : (8'hb4))) ?
                  $signed(wire652[(1'h1):(1'h0)]) : (~&($signed(wire276[(4'hc):(2'h2)]) * $unsigned((|wire668)))));
            end
          if ($signed((8'hb4)))
            begin
              reg674 <= $signed(reg671[(1'h1):(1'h1)]);
              reg675 <= reg672;
              reg676 <= ((~|reg674) ?
                  (wire652[(3'h6):(1'h0)] ~^ $signed($unsigned(reg673))) : ($signed((&(reg661 >>> wire275))) ?
                      $signed((wire275[(4'h8):(1'h1)] ?
                          $unsigned(wire652) : {wire652})) : wire276[(4'hb):(3'h4)]));
              reg677 = $unsigned($unsigned(({{reg671,
                      wire275}} ^~ (~wire275[(3'h6):(1'h1)]))));
            end
          else
            begin
              reg674 <= {$unsigned((wire652[(4'h8):(3'h7)] ?
                      reg663[(3'h5):(1'h1)] : $signed((wire275 - wire653))))};
              reg677 = (reg663 ? $signed((8'h9c)) : $unsigned(wire650));
              reg678 <= {$signed({{reg670[(4'hf):(4'hd)]},
                      reg670[(1'h0):(1'h0)]})};
              reg679 <= (wire274[(3'h7):(3'h7)] ?
                  (((+$signed(forvar669)) || $unsigned((wire668 ?
                          (8'haa) : reg673))) ?
                      $unsigned((wire274 + reg667[(4'hf):(4'h9)])) : ((^~$signed((8'hbd))) ?
                          {$unsigned(reg658)} : ($signed(reg658) ?
                              forvar669 : wire277))) : $signed({reg673,
                      (~^wire275)}));
              reg680 = ({($signed($unsigned((7'h40))) ?
                          wire277[(4'hd):(4'ha)] : (reg673[(5'h10):(4'h9)] ~^ (reg666 ?
                              reg673 : wire650))),
                      (($signed(reg658) * (~wire275)) ?
                          wire276 : $signed($unsigned(reg666)))} ?
                  $unsigned((~&(reg663[(2'h3):(1'h0)] ~^ {reg675}))) : (|(&{$signed(reg663),
                      (wire650 < wire276)})));
            end
          reg681 = (reg679[(4'hd):(4'hd)] ? reg663 : wire277);
        end
      for (forvar682 = (1'h0); (forvar682 < (1'h1)); forvar682 = (forvar682 + (1'h1)))
        begin
          if ({forvar682})
            begin
              reg683 <= forvar682;
              reg684 <= $unsigned($unsigned((8'hab)));
              reg685 <= wire668;
            end
          else
            begin
              reg686 = (|reg678[(3'h6):(3'h6)]);
            end
          reg687 = $signed($signed(((reg671 ?
                  (wire276 ? reg667 : wire277) : (forvar682 ?
                      wire668 : reg670)) ?
              {wire276[(3'h6):(1'h1)], reg673} : (~|(wire278 - reg678)))));
        end
      for (forvar688 = (1'h0); (forvar688 < (2'h3)); forvar688 = (forvar688 + (1'h1)))
        begin
          reg689 = (reg666[(3'h4):(2'h2)] | reg687);
          if ($signed(({((reg674 ? wire277 : reg679) ?
                      $signed(reg683) : {(8'hbd), wire668})} ?
              (~&(+reg670[(5'h11):(2'h2)])) : reg675)))
            begin
              reg690 = wire275[(2'h3):(1'h1)];
            end
          else
            begin
              reg691 <= $unsigned($signed((^~(~|(wire277 ?
                  (8'hb9) : reg679)))));
              reg692 <= ((reg667 < $unsigned($unsigned($unsigned(wire652)))) > wire276[(4'h8):(2'h2)]);
              reg693 <= (|((8'h9c) ?
                  $unsigned((~(reg678 >= wire277))) : ((~&$unsigned(reg691)) ?
                      $unsigned(reg658) : (reg683[(3'h4):(2'h2)] && (~^reg675)))));
            end
          reg694 = ((|$signed(((reg663 == wire668) ?
                  (wire274 ? wire276 : reg680) : (wire668 ?
                      reg680 : reg658)))) ?
              $unsigned((reg690[(3'h6):(1'h0)] ?
                  reg672 : forvar669)) : reg693[(3'h6):(1'h1)]);
          reg695 <= {reg661,
              ((!((8'ha1) > {wire650})) ?
                  {(((7'h43) >= wire652) && (reg672 * reg671))} : {wire652[(3'h6):(2'h2)],
                      ($signed(reg691) ?
                          (reg692 ~^ (8'hab)) : $unsigned(reg677))})};
          if (({$unsigned($signed(reg661[(3'h4):(2'h2)])),
                  (^~$unsigned((~^reg673)))} ?
              wire276[(1'h0):(1'h0)] : (|(~^(|((7'h49) <<< reg691))))))
            begin
              reg696 = wire668;
            end
          else
            begin
              reg697 <= $signed(($unsigned(reg695[(2'h2):(1'h0)]) ?
                  (-(reg672 << (reg666 | reg696))) : $unsigned($signed(((8'hb8) <<< reg680)))));
              reg698 = (-(8'ha8));
              reg699 <= (8'hbb);
              reg700 = ($unsigned((8'haa)) >> (^~($unsigned(reg696) >= (reg687 ?
                  (reg690 ? reg666 : reg670) : (wire277 ? reg693 : reg667)))));
              reg701 = reg674[(1'h0):(1'h0)];
            end
        end
      reg702 <= $unsigned((reg696 ?
          $unsigned(reg661[(2'h3):(1'h1)]) : {reg666[(1'h0):(1'h0)]}));
    end
  module703 #() modinst1316 (wire1315, clk, reg667, reg678, wire668, reg674, reg695);
  module1025 #() modinst1318 (.wire1028(reg684), .clk(clk), .wire1029(reg674), .wire1027(reg675), .wire1026(reg679), .y(wire1317), .wire1030(reg658));
  always
    @(posedge clk) begin
      reg1319 <= reg679[(4'he):(4'h9)];
      reg1320 = {$unsigned(wire274[(1'h1):(1'h0)]),
          (reg674 ?
              $unsigned(((8'hb9) ?
                  reg663[(2'h3):(1'h0)] : {reg691})) : (reg658 ?
                  $unsigned((reg691 + (8'hac))) : {reg675[(4'ha):(4'h8)],
                      wire668}))};
      reg1321 = (!wire278[(3'h6):(2'h2)]);
      for (forvar1322 = (1'h0); (forvar1322 < (2'h2)); forvar1322 = (forvar1322 + (1'h1)))
        begin
          reg1323 <= ((reg671 < (reg671[(5'h10):(2'h2)] >= ($signed(reg675) <<< (reg1319 == reg663)))) + ((reg674 ~^ (8'haf)) < wire275[(5'h11):(4'h9)]));
          for (forvar1324 = (1'h0); (forvar1324 < (2'h3)); forvar1324 = (forvar1324 + (1'h1)))
            begin
              reg1325 <= (!{reg691[(3'h5):(3'h4)]});
              reg1326 = $signed($signed((^~$signed((+(7'h4a))))));
              reg1327 <= {wire277[(2'h2):(1'h0)]};
            end
          reg1328 = reg1320[(1'h0):(1'h0)];
          reg1329 <= reg1320[(1'h1):(1'h0)];
        end
      reg1330 <= $signed(reg667);
    end
  always
    @(posedge clk) begin
      if ((8'had))
        begin
          if ((7'h49))
            begin
              reg1331 <= {$signed(((wire274 ?
                          (reg1319 ? wire1317 : (8'hab)) : reg685) ?
                      (reg1330 ?
                          (reg676 >> wire668) : $signed(reg678)) : reg1319)),
                  (((&$unsigned(reg1330)) ?
                      (!wire652[(1'h0):(1'h0)]) : (!reg674)) && (wire278[(5'h11):(4'hd)] ?
                      $signed((reg693 <<< wire278)) : (~|(-(7'h47)))))};
              reg1332 = (reg667[(5'h12):(3'h5)] <<< (reg670 ?
                  $unsigned($signed(wire1315[(4'hf):(4'h8)])) : (~^$signed(reg1325[(4'h9):(2'h3)]))));
              reg1333 <= $signed(reg695);
              reg1334 <= ($unsigned((((reg1333 ?
                  wire653 : reg679) * reg676[(5'h15):(5'h15)]) >= $unsigned((reg683 & wire276)))) < $unsigned((reg695[(4'hf):(4'hc)] ~^ wire274)));
            end
          else
            begin
              reg1331 <= ($unsigned((((wire1315 ?
                      wire1317 : reg684) <= {(8'hb9)}) ?
                  ({(8'hbf),
                      reg693} * $unsigned(reg679)) : (wire1317[(3'h4):(2'h3)] ?
                      reg1323[(3'h7):(3'h7)] : reg1330[(5'h14):(3'h6)]))) > ((~$signed({reg661})) < $unsigned(reg679)));
              reg1332 = (reg667 >= (~reg685));
              reg1333 <= (!((($signed((7'h4a)) ?
                          (reg1331 ? reg1334 : wire668) : reg693) ?
                      (((8'h9e) ? (8'hbc) : (8'h9f)) ?
                          (reg695 && wire274) : reg661[(1'h1):(1'h1)]) : ($unsigned(wire650) ?
                          {reg658} : $unsigned(reg692))) ?
                  {(reg695[(4'h9):(2'h2)] ? wire1317 : (reg1332 ~^ reg699)),
                      wire276[(4'hd):(4'h8)]} : ((^~$signed(reg1329)) ?
                      $signed($signed(reg1332)) : ((reg691 || reg685) ?
                          (~&reg661) : (reg683 <= reg683)))));
              reg1334 <= reg1325;
            end
          reg1335 <= $signed(reg692);
          reg1336 = wire1315;
        end
      else
        begin
          if ({reg1336})
            begin
              reg1332 = $unsigned(((((^~reg676) ?
                      (-reg663) : $unsigned(wire1317)) <<< reg661[(3'h4):(2'h2)]) ?
                  reg1327 : (^~$signed((wire1317 || (7'h49))))));
              reg1333 <= (wire274 | ((^~reg702) + $signed((~|(reg663 ?
                  (8'hb7) : reg679)))));
              reg1336 = (~^reg683);
            end
          else
            begin
              reg1331 <= (~&{($signed($signed(wire274)) ?
                      reg670[(1'h1):(1'h0)] : (reg675 << $signed(reg1329))),
                  (^~reg1333[(4'ha):(4'h9)])});
            end
          for (forvar1337 = (1'h0); (forvar1337 < (1'h1)); forvar1337 = (forvar1337 + (1'h1)))
            begin
              reg1338 <= (8'hbe);
              reg1339 <= reg1336[(3'h7):(3'h7)];
              reg1340 <= $signed((|(&$unsigned(reg685))));
            end
          for (forvar1341 = (1'h0); (forvar1341 < (1'h0)); forvar1341 = (forvar1341 + (1'h1)))
            begin
              reg1342 <= (|$unsigned((7'h48)));
              reg1343 <= $unsigned($unsigned((reg695[(4'ha):(4'h9)] ^ (wire652[(4'h8):(1'h1)] < reg1329))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg1344 = $signed(reg1327[(3'h5):(3'h5)]);
    end
  assign wire1345 = wire650[(5'h18):(5'h12)];
  assign wire1346 = ($signed(($signed($signed((7'h42))) || ((8'hab) ?
                            reg692 : $unsigned(reg702)))) ?
                        $unsigned(((~^(wire276 ? (8'hae) : reg678)) ?
                            $unsigned((8'hac)) : (-(wire652 || wire278)))) : (&$signed((wire275[(5'h11):(1'h0)] ?
                            (7'h47) : reg1323))));
  always
    @(posedge clk) begin
      reg1347 <= reg1334;
      if (reg675)
        begin
          if ((8'hba))
            begin
              reg1348 <= (!reg1330[(4'hc):(3'h4)]);
            end
          else
            begin
              reg1348 <= reg1335;
              reg1349 <= ($unsigned((wire668[(4'hb):(4'h8)] ?
                      ((reg699 <= reg1342) ?
                          (~^(7'h49)) : $unsigned(wire274)) : reg1330[(4'hb):(4'hb)])) ?
                  $signed(($unsigned($signed(reg1335)) ?
                      {reg1329, wire277[(4'hf):(1'h1)]} : {reg1338,
                          (!(8'had))})) : wire1317[(4'hd):(4'h8)]);
              reg1350 <= ($signed({wire274[(4'hc):(2'h2)],
                  (wire1315[(5'h12):(4'hd)] ?
                      {(7'h45)} : $unsigned(reg676))}) <= $signed((^~wire275)));
              reg1351 = $signed($unsigned($signed(((wire1346 << wire653) >>> (|reg1325)))));
            end
          if (((wire1346[(3'h5):(3'h4)] ?
                  ({(8'ha0)} || $signed({wire275, reg674})) : ((&(+wire1345)) ?
                      $unsigned($signed(wire274)) : ($unsigned(reg670) & (reg1342 ?
                          reg1331 : reg666)))) ?
              $unsigned($unsigned((!(reg1342 | reg699)))) : wire1346[(1'h0):(1'h0)]))
            begin
              reg1352 <= $signed((!reg1340));
            end
          else
            begin
              reg1353 = $signed((wire1315 >= $unsigned(reg1338)));
              reg1354 = reg670[(3'h4):(1'h0)];
              reg1355 <= $unsigned((~&(reg1349 ^ (~&$unsigned((8'h9c))))));
            end
          reg1356 = reg683;
        end
      else
        begin
          reg1348 <= $signed(reg1329[(4'hb):(4'hb)]);
          reg1351 = ($signed(({(-(8'ha3)), (reg671 ? reg1334 : (8'ha4))} ?
                  $unsigned((reg1327 & reg1339)) : {$signed(reg658),
                      (~reg1335)})) ?
              (reg1356 ~^ ((&(~^(8'ha3))) ?
                  $signed((^~reg1330)) : $unsigned(((8'ha7) ?
                      reg674 : reg667)))) : reg675);
          reg1352 <= $signed((($signed(reg1319[(1'h0):(1'h0)]) ^ $signed((wire1317 ?
                  reg692 : wire274))) ?
              reg1348[(4'h9):(4'h9)] : wire652[(3'h5):(1'h0)]));
          for (forvar1353 = (1'h0); (forvar1353 < (1'h1)); forvar1353 = (forvar1353 + (1'h1)))
            begin
              reg1355 <= $unsigned((8'haf));
              reg1357 <= $unsigned((~^(^~(8'hbf))));
              reg1358 = ((~|$signed((7'h44))) ^ ((|($unsigned(reg684) && (reg1327 ?
                  reg1327 : (7'h42)))) >= $signed(($unsigned(reg674) ?
                  reg1334 : $signed(reg1349)))));
              reg1359 = wire653;
            end
        end
    end
  always
    @(posedge clk) begin
      reg1360 <= $signed(reg1357);
      for (forvar1361 = (1'h0); (forvar1361 < (1'h0)); forvar1361 = (forvar1361 + (1'h1)))
        begin
          for (forvar1362 = (1'h0); (forvar1362 < (3'h4)); forvar1362 = (forvar1362 + (1'h1)))
            begin
              reg1363 <= (-$signed($signed(wire668[(5'h10):(5'h10)])));
              reg1364 = $unsigned((7'h42));
              reg1365 <= ((({$signed((7'h48)),
                      $unsigned(reg1349)} != $signed((reg1342 ?
                      reg678 : reg695))) & (~reg1347[(4'hc):(1'h1)])) ?
                  ({reg1364[(3'h7):(3'h4)], (~|wire1315)} > ((reg658 ?
                          (^(7'h41)) : (reg678 ? reg702 : (7'h45))) ?
                      $unsigned(reg1319[(2'h3):(2'h3)]) : (wire275 << (reg1343 ^~ forvar1361)))) : (!(^(reg1364[(1'h0):(1'h0)] != reg667[(5'h10):(3'h7)]))));
            end
          if ($signed(reg670))
            begin
              reg1366 <= {(((reg1334[(4'ha):(2'h2)] != {reg1365}) >>> reg1349) && $unsigned(reg670))};
              reg1367 <= $unsigned((reg1350 && {$signed((|(7'h47))),
                  (|{reg1347, reg1350})}));
              reg1368 = (wire653 ? wire274 : reg1327);
              reg1369 <= (~reg693);
            end
          else
            begin
              reg1366 <= (reg1364[(2'h2):(2'h2)] ^ $signed(reg1357[(3'h5):(2'h3)]));
            end
          reg1370 <= reg1369[(3'h6):(3'h5)];
        end
      reg1371 = reg1366;
    end
  always
    @(posedge clk) begin
      reg1372 <= (-$unsigned(($signed((reg1350 == reg1355)) ?
          (8'hb1) : ((reg1369 || wire1315) == $unsigned(wire275)))));
      reg1373 <= ({(~(reg692 ? {(8'haa)} : (+reg1365)))} ?
          $signed($unsigned($signed(reg1347[(3'h4):(2'h2)]))) : $unsigned(reg684[(2'h3):(2'h2)]));
      if ((-(^$signed(((reg658 ? (7'h43) : reg658) >= (~^reg1333))))))
        begin
          reg1374 <= ({reg697} ~^ {((^$unsigned(reg1333)) <= {{reg679, reg1349},
                  reg1367})});
          if (reg1369[(3'h6):(3'h4)])
            begin
              reg1375 = (reg661 <= $unsigned($unsigned((&$unsigned(wire274)))));
              reg1376 = $unsigned(($unsigned($signed((reg1367 || reg1335))) ^ $signed((~^(reg661 != wire653)))));
            end
          else
            begin
              reg1377 <= $unsigned((((reg1370[(4'hb):(3'h6)] ?
                      (reg1319 && reg1327) : (~reg1334)) ?
                  reg1357 : reg1360) * $signed(reg671[(4'hf):(4'ha)])));
            end
          for (forvar1378 = (1'h0); (forvar1378 < (1'h0)); forvar1378 = (forvar1378 + (1'h1)))
            begin
              reg1379 = (+{$unsigned(((~|reg1352) + $signed(reg695))),
                  ((-(+wire275)) ?
                      $signed($signed(wire650)) : wire274[(4'h8):(4'h8)])});
              reg1380 = $unsigned({(+((reg1376 ^~ wire668) ?
                      (reg1333 >> reg1342) : reg1377[(2'h2):(1'h1)])),
                  (($signed((8'hbc)) ^~ (reg1374 >= reg674)) | $signed((-reg693)))});
            end
        end
      else
        begin
          if ((reg693 == {reg1360}))
            begin
              reg1375 = reg692[(3'h4):(1'h0)];
              reg1377 <= $signed(reg1366);
            end
          else
            begin
              reg1375 = ((($signed(reg1330) ?
                  reg1325[(5'h10):(2'h3)] : $signed($unsigned(reg1369))) ^ reg697[(3'h5):(1'h0)]) >>> (($signed(reg1333) >>> ({wire277} ?
                  reg1333 : $unsigned(reg1323))) <= (($unsigned((8'ha6)) - $signed(reg1376)) ?
                  ({reg1339} + (reg676 ? wire275 : (8'ha1))) : reg1376)));
              reg1377 <= reg1357;
            end
          if ({$signed(reg1339[(3'h4):(1'h1)]),
              $signed(({(reg663 ^~ reg1334)} ?
                  $signed($unsigned(reg1335)) : (8'ha6)))})
            begin
              reg1378 <= ((^reg661) ?
                  {(reg1331 > ((reg1340 ? reg1335 : reg1350) >>> (|reg1333))),
                      ($unsigned((wire1345 ?
                          reg679 : reg658)) != ($signed(reg1370) != (reg1380 ?
                          reg1370 : reg1377)))} : ({reg1333[(1'h0):(1'h0)],
                          (((8'hb8) - (8'ha0)) <<< {reg684})} ?
                      $signed(reg1357) : $signed((8'hb3))));
              reg1379 = (reg683[(1'h0):(1'h0)] ?
                  (!$signed(reg1379)) : ((-wire277) ?
                      {$signed({reg1372}),
                          $unsigned(reg691[(4'h8):(3'h7)])} : {$unsigned((8'hb7)),
                          $signed(reg1355[(3'h5):(2'h2)])}));
              reg1381 <= (8'haf);
              reg1382 = (reg1338 ^ ((!$unsigned($signed(reg692))) ?
                  reg1370[(4'h9):(4'h9)] : reg695[(4'hf):(2'h3)]));
              reg1383 <= reg679[(3'h7):(2'h2)];
            end
          else
            begin
              reg1378 <= ((wire653[(3'h6):(2'h3)] ?
                      (^~((reg658 & reg1360) >= (8'hb7))) : $signed({(~&reg693)})) ?
                  reg1372 : (8'ha4));
              reg1379 = $unsigned((+(!$unsigned($unsigned(reg1369)))));
              reg1381 <= reg699;
              reg1382 = (~^$signed((~&(^reg1379[(3'h7):(1'h1)]))));
              reg1384 = {reg1378};
            end
          for (forvar1385 = (1'h0); (forvar1385 < (3'h4)); forvar1385 = (forvar1385 + (1'h1)))
            begin
              reg1386 <= ($unsigned(reg1380) ? reg702 : $signed(wire1345));
              reg1387 <= $signed((($unsigned($signed(reg1369)) || $signed(reg1333[(4'ha):(1'h1)])) >> (8'hac)));
            end
          for (forvar1388 = (1'h0); (forvar1388 < (1'h0)); forvar1388 = (forvar1388 + (1'h1)))
            begin
              reg1389 = reg671;
              reg1390 = (reg674[(5'h14):(3'h5)] ^ wire275);
              reg1391 = $signed($signed((forvar1388 && reg678)));
              reg1392 = reg1325[(5'h12):(2'h2)];
              reg1393 <= $signed(((reg1323[(2'h2):(1'h0)] ?
                      $signed((~wire652)) : $unsigned((forvar1385 ?
                          reg699 : reg675))) ?
                  (~^$unsigned({reg1330})) : (((~|reg1369) >>> reg683[(3'h7):(2'h3)]) && $unsigned(reg658[(3'h4):(3'h4)]))));
            end
          if ((+$unsigned(reg1335[(4'he):(4'h9)])))
            begin
              reg1394 = reg1343;
              reg1395 <= (~|$unsigned($signed($signed((reg1372 || reg1327)))));
              reg1396 <= reg1329[(3'h5):(1'h1)];
              reg1397 = {(({reg692, $signed(reg1381)} ?
                          wire1315 : ($unsigned(reg695) > (8'hb7))) ?
                      {{wire276[(3'h4):(2'h2)]},
                          reg1333[(1'h0):(1'h0)]} : {{((8'ha2) >= reg1339)}})};
              reg1398 = (~|(reg679 > wire276[(4'h8):(1'h0)]));
            end
          else
            begin
              reg1395 <= (&reg1333);
              reg1397 = $signed(reg1378[(4'hc):(3'h5)]);
              reg1399 <= {(8'h9e)};
            end
        end
      for (forvar1400 = (1'h0); (forvar1400 < (1'h1)); forvar1400 = (forvar1400 + (1'h1)))
        begin
          reg1401 = (reg1375[(4'hf):(4'h9)] == $signed(reg1391[(2'h2):(1'h1)]));
        end
      for (forvar1402 = (1'h0); (forvar1402 < (2'h2)); forvar1402 = (forvar1402 + (1'h1)))
        begin
          for (forvar1403 = (1'h0); (forvar1403 < (3'h4)); forvar1403 = (forvar1403 + (1'h1)))
            begin
              reg1404 <= (8'hab);
              reg1405 <= reg1366;
              reg1406 = ((~$signed($signed($unsigned(forvar1403)))) ?
                  wire278[(3'h4):(2'h3)] : ((~(reg1391 >= (reg676 ?
                          forvar1385 : reg1382))) ?
                      (8'hb6) : (forvar1385[(1'h1):(1'h1)] != reg1398[(3'h7):(3'h5)])));
              reg1407 <= (^(reg679[(1'h0):(1'h0)] <= reg1327));
              reg1408 <= $unsigned(reg684);
            end
        end
    end
  module279 #() modinst1410 (.wire283(reg1377), .wire282(wire652), .wire284(reg1352), .wire281(reg699), .y(wire1409), .wire280(reg1404), .clk(clk));
  module1192 #() modinst1412 (wire1411, clk, reg1327, reg670, reg1367, reg658, reg1387);
  always
    @(posedge clk) begin
      reg1413 = $signed($signed((~&{(reg675 > reg1381)})));
      for (forvar1414 = (1'h0); (forvar1414 < (2'h3)); forvar1414 = (forvar1414 + (1'h1)))
        begin
          if ((reg1399 >= (+(&$signed(((8'ha5) ? reg1319 : (7'h4a)))))))
            begin
              reg1415 <= $unsigned(reg1404);
              reg1416 <= $unsigned($signed($unsigned(reg1405)));
              reg1417 <= $signed(wire1409[(3'h5):(1'h1)]);
              reg1418 = $signed({reg676});
              reg1419 = ($unsigned((^~wire650)) ?
                  {$unsigned($signed((reg1377 ^ reg1366)))} : ((+$signed($unsigned((8'ha1)))) < {$signed($signed(reg1334))}));
            end
          else
            begin
              reg1415 <= (reg1365[(1'h1):(1'h1)] ?
                  reg1329[(1'h1):(1'h0)] : (reg663 ?
                      reg658 : (((reg1325 ? reg695 : wire1411) ?
                              {reg1360, reg1419} : $unsigned(reg1405)) ?
                          ((reg1333 ? (8'ha3) : wire276) ?
                              $signed((8'hbb)) : (reg678 ?
                                  reg1387 : reg1339)) : reg1340)));
              reg1418 = {(+wire1317[(5'h14):(5'h12)])};
            end
          if ((reg1413[(3'h5):(2'h3)] ?
              $signed((|(wire1345 >>> reg1333))) : ((reg679[(4'hc):(3'h4)] || {{wire653,
                      reg1417}}) ~^ $unsigned(wire668[(4'hf):(3'h4)]))))
            begin
              reg1420 <= {reg1386};
              reg1421 <= reg671[(4'hc):(4'ha)];
              reg1422 <= reg1325[(4'he):(4'ha)];
              reg1423 <= (!$signed(reg1365[(3'h5):(3'h4)]));
              reg1424 <= reg1418[(3'h7):(2'h2)];
            end
          else
            begin
              reg1425 = $signed($unsigned($signed((8'ha3))));
              reg1426 = ((8'ha4) ? (8'hb0) : reg1335);
              reg1427 = (($unsigned(((^reg1413) - reg1417)) >>> reg674[(5'h12):(4'hb)]) ?
                  ({{reg1387, reg693}} ?
                      $signed(reg1415) : (~^$signed($unsigned(reg1405)))) : (reg663[(3'h5):(2'h3)] || {((reg1413 != (8'hb5)) & {reg1404})}));
              reg1428 <= {($signed((reg1395[(2'h2):(1'h1)] ?
                      $unsigned(reg693) : {reg1419})) - reg1377)};
              reg1429 = reg670;
            end
          for (forvar1430 = (1'h0); (forvar1430 < (2'h3)); forvar1430 = (forvar1430 + (1'h1)))
            begin
              reg1431 <= (reg670 ?
                  ($unsigned((~{reg1428})) <<< wire1317[(5'h13):(5'h10)]) : (!{({reg1372} ?
                          reg702 : reg683[(3'h4):(2'h3)])}));
            end
          if ((8'hac))
            begin
              reg1432 = $signed($unsigned(($unsigned((wire650 ?
                      reg1381 : (8'ha8))) ?
                  reg1407[(4'hb):(4'hb)] : reg1323[(4'hd):(3'h4)])));
              reg1433 <= reg1319;
              reg1434 <= $unsigned((~|($unsigned($unsigned(reg1350)) << $signed($unsigned((7'h49))))));
              reg1435 <= $signed(reg1421[(3'h4):(1'h0)]);
              reg1436 = ((^($signed((reg1399 >= reg1360)) & $unsigned((wire650 ^~ reg1367)))) * $signed(reg1365));
            end
          else
            begin
              reg1433 <= $unsigned(((reg666[(1'h1):(1'h0)] >> (reg699 ?
                  $unsigned(reg1419) : (reg1378 >> reg671))) & $signed($signed((|reg658)))));
              reg1434 <= reg699;
              reg1435 <= ({$signed(((!(7'h44)) > (~&(8'hb6)))),
                  wire275} || (((~&(reg661 ? reg1418 : reg1355)) ?
                      (+(reg1365 ? reg685 : reg666)) : wire652[(3'h6):(1'h1)]) ?
                  $signed(((reg1431 >= reg1435) * (reg1330 ?
                      reg1425 : wire278))) : (^((-reg1357) <= reg685[(2'h3):(2'h3)]))));
              reg1437 <= reg678[(2'h3):(1'h0)];
            end
          if (reg1335[(4'h8):(3'h7)])
            begin
              reg1438 <= wire276[(4'h9):(2'h3)];
              reg1439 = reg661;
              reg1440 = (wire1345 ?
                  ((~|(~&reg691)) >> $unsigned((reg675[(2'h2):(1'h1)] ^~ $unsigned(reg1383)))) : (~|$unsigned({(reg1439 != reg1428)})));
              reg1441 = ($signed(($signed(reg1433) ?
                      (|$signed(reg1415)) : reg666)) ?
                  ($signed(((wire668 == reg1404) ^~ wire650)) >= {$signed(reg1350[(2'h2):(1'h1)])}) : $unsigned($unsigned($unsigned(wire650))));
              reg1442 <= reg1429;
            end
          else
            begin
              reg1439 = (($signed(wire1317[(5'h14):(4'hb)]) ^ (($signed(reg685) >>> (-reg676)) ^ (~(reg1350 | reg1378)))) ?
                  $unsigned({((reg667 ? reg1338 : (8'ha3)) ?
                          reg1329 : $unsigned(reg685)),
                      ((~^reg1339) + $signed(reg1386))}) : {(~^reg1439[(4'ha):(3'h5)])});
              reg1440 = $unsigned(($signed($signed((reg1363 << reg1442))) > ((^(reg1349 ?
                  reg1333 : reg1330)) || $unsigned(reg1343))));
              reg1441 = (reg1419 ?
                  (reg1365[(3'h4):(2'h3)] == reg1334) : $unsigned((~^$signed((!reg1319)))));
            end
        end
      for (forvar1443 = (1'h0); (forvar1443 < (3'h4)); forvar1443 = (forvar1443 + (1'h1)))
        begin
          reg1444 <= $signed({$unsigned((&(|reg1439))),
              $unsigned({$unsigned(wire653), reg1419[(4'h8):(3'h5)]})});
          for (forvar1445 = (1'h0); (forvar1445 < (2'h3)); forvar1445 = (forvar1445 + (1'h1)))
            begin
              reg1446 <= (~$signed($unsigned($unsigned((&(7'h46))))));
              reg1447 = $signed((^~$unsigned($unsigned((~^reg1331)))));
            end
          for (forvar1448 = (1'h0); (forvar1448 < (1'h0)); forvar1448 = (forvar1448 + (1'h1)))
            begin
              reg1449 <= (|((($unsigned(forvar1448) & reg675) >= $signed($signed(reg1415))) >>> (8'hb4)));
              reg1450 = (~|(({reg1339[(3'h4):(3'h4)]} ^ (8'ha5)) - {(~&(reg1327 ?
                      reg1396 : reg1374))}));
            end
        end
      reg1451 <= ($unsigned(($unsigned(reg1432) ?
          reg1329 : forvar1445)) <<< wire650);
      reg1452 = reg1439[(3'h6):(3'h4)];
    end
  module1025 #() modinst1454 (.wire1029(reg1363), .wire1030(reg1355), .wire1027(reg1435), .wire1026(reg1331), .y(wire1453), .wire1028(reg1334), .clk(clk));
  always
    @(posedge clk) begin
      reg1455 <= ({reg666,
          (reg1428[(5'h12):(1'h0)] ?
              $unsigned(reg1383[(1'h0):(1'h0)]) : $unsigned($signed((8'hb7))))} ^ (8'hba));
      for (forvar1456 = (1'h0); (forvar1456 < (1'h1)); forvar1456 = (forvar1456 + (1'h1)))
        begin
          reg1457 <= $signed(reg1417);
          if (reg1435)
            begin
              reg1458 <= (8'haf);
              reg1459 = (reg1327[(5'h14):(5'h12)] ?
                  $unsigned($unsigned(((reg1323 ? reg1374 : reg1444) ?
                      reg1378 : $unsigned((7'h42))))) : $signed($unsigned(((reg1373 | reg697) ?
                      reg1357[(3'h4):(3'h4)] : (reg1437 ?
                          reg1323 : (7'h47))))));
            end
          else
            begin
              reg1459 = (reg1329[(4'hf):(4'hf)] ^ $unsigned((reg1350 ?
                  (((8'hb6) ? reg1335 : reg1433) ?
                      (reg1446 - reg1325) : $signed(reg1363)) : ((~&reg1395) ?
                      reg692 : ((8'hbb) ? reg1369 : reg1366)))));
              reg1460 <= {reg1343,
                  (($unsigned((reg1323 - reg1349)) ?
                      $unsigned(reg1350) : ({wire1317, reg1338} ?
                          reg1408[(2'h3):(2'h3)] : {reg1393,
                              (8'ha1)})) ^~ reg667)};
            end
          reg1461 <= reg679[(1'h1):(1'h1)];
          for (forvar1462 = (1'h0); (forvar1462 < (2'h3)); forvar1462 = (forvar1462 + (1'h1)))
            begin
              reg1463 <= reg1431;
              reg1464 <= ($unsigned($unsigned(reg1327)) | ((((-reg1408) != $signed(reg1334)) ?
                  wire652 : {$unsigned(reg1395)}) == reg1335));
            end
          reg1465 = $unsigned($unsigned((({reg1367, reg1370} ?
                  (-reg667) : $signed(wire275)) ?
              (&(wire1317 > reg1352)) : (^~reg1442[(5'h16):(3'h4)]))));
        end
      reg1466 = $signed(forvar1456);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module703
#(parameter param1313 = ({(~|({(7'h40)} ? {(8'haa)} : (!(8'hbf))))} ? (~&(|{{(8'ha8), (8'hbd)}, (^~(7'h44))})) : (~&(8'ha6))), 
parameter param1314 = (((^(param1313 >= (param1313 ? param1313 : param1313))) ? {((param1313 - param1313) ? (param1313 ? param1313 : param1313) : ((8'hb6) >> param1313))} : {(param1313 ? {param1313, param1313} : param1313)}) ? ((~|(-(8'hb4))) ? (param1313 <<< param1313) : (|param1313)) : (((param1313 ? param1313 : (^param1313)) ? {param1313, ((8'hb3) ? param1313 : (7'h41))} : (+{(8'hb6), (7'h40)})) ? (((param1313 << (8'hba)) ^ (param1313 >> param1313)) ? ((^~param1313) ? ((8'ha1) ? (8'h9f) : param1313) : (param1313 - (8'hb5))) : ((param1313 ? param1313 : param1313) >> {param1313})) : (((|param1313) >> ((7'h4a) ? param1313 : param1313)) - (param1313 ? (param1313 & param1313) : {param1313, param1313})))))
(y, clk, wire704, wire705, wire706, wire707, wire708);
  output wire [(32'h68a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire704;
  input wire signed [(5'h16):(1'h0)] wire705;
  input wire [(5'h17):(1'h0)] wire706;
  input wire [(5'h11):(1'h0)] wire707;
  input wire [(4'hf):(1'h0)] wire708;
  wire [(5'h11):(1'h0)] wire1312;
  wire [(3'h4):(1'h0)] wire1167;
  wire [(2'h2):(1'h0)] wire821;
  wire signed [(5'h12):(1'h0)] wire823;
  wire signed [(4'h9):(1'h0)] wire824;
  wire [(3'h7):(1'h0)] wire825;
  wire signed [(5'h12):(1'h0)] wire862;
  wire [(4'h9):(1'h0)] wire994;
  wire signed [(4'hb):(1'h0)] wire1169;
  wire [(5'h12):(1'h0)] wire1170;
  wire [(5'h13):(1'h0)] wire1171;
  wire [(5'h16):(1'h0)] wire1190;
  wire signed [(5'h11):(1'h0)] wire1191;
  wire [(3'h5):(1'h0)] wire1288;
  wire [(5'h15):(1'h0)] wire1290;
  wire signed [(5'h10):(1'h0)] wire1292;
  reg [(4'h8):(1'h0)] reg1311 = (1'h0);
  reg [(5'h15):(1'h0)] reg1310 = (1'h0);
  reg [(4'h9):(1'h0)] reg1308 = (1'h0);
  reg [(4'hd):(1'h0)] reg1307 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1304 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1303 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1300 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1299 = (1'h0);
  reg [(5'h17):(1'h0)] reg1296 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1187 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1186 = (1'h0);
  reg [(5'h17):(1'h0)] reg1185 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1179 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1183 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1177 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1175 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1174 = (1'h0);
  reg [(3'h4):(1'h0)] reg1172 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1020 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1019 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1017 = (1'h0);
  reg [(5'h18):(1'h0)] reg1014 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1011 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1010 = (1'h0);
  reg [(4'h9):(1'h0)] reg1008 = (1'h0);
  reg [(3'h7):(1'h0)] reg1007 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1005 = (1'h0);
  reg [(4'hd):(1'h0)] reg1003 = (1'h0);
  reg [(5'h15):(1'h0)] reg999 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg998 = (1'h0);
  reg [(4'hc):(1'h0)] reg826 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg827 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg829 = (1'h0);
  reg [(5'h17):(1'h0)] reg831 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg832 = (1'h0);
  reg [(4'h9):(1'h0)] reg837 = (1'h0);
  reg [(5'h10):(1'h0)] reg838 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg839 = (1'h0);
  reg [(4'h8):(1'h0)] reg841 = (1'h0);
  reg signed [(4'he):(1'h0)] reg846 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg848 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg851 = (1'h0);
  reg [(5'h13):(1'h0)] reg852 = (1'h0);
  reg [(4'ha):(1'h0)] reg854 = (1'h0);
  reg [(5'h15):(1'h0)] reg857 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg858 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg859 = (1'h0);
  reg [(5'h11):(1'h0)] reg861 = (1'h0);
  reg [(5'h16):(1'h0)] reg1309 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1306 = (1'h0);
  reg [(4'he):(1'h0)] reg1305 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1302 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1301 = (1'h0);
  reg [(5'h12):(1'h0)] reg1298 = (1'h0);
  reg [(3'h4):(1'h0)] reg1297 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1295 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1294 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1189 = (1'h0);
  reg [(4'hb):(1'h0)] reg1188 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1184 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1182 = (1'h0);
  reg [(4'hf):(1'h0)] reg1181 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1180 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1179 = (1'h0);
  reg [(4'h9):(1'h0)] reg1178 = (1'h0);
  reg [(5'h17):(1'h0)] reg1176 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1173 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1024 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1023 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1022 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1021 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1018 = (1'h0);
  reg [(4'he):(1'h0)] reg1016 = (1'h0);
  reg [(4'h8):(1'h0)] reg1015 = (1'h0);
  reg [(4'hc):(1'h0)] reg1013 = (1'h0);
  reg [(4'he):(1'h0)] reg1012 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1009 = (1'h0);
  reg [(5'h10):(1'h0)] reg1006 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1004 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1002 = (1'h0);
  reg [(5'h17):(1'h0)] reg1001 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1000 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar997 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg996 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg860 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg856 = (1'h0);
  reg [(4'hd):(1'h0)] reg855 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar853 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg850 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg849 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar847 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg845 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg844 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg833 = (1'h0);
  reg [(5'h10):(1'h0)] forvar826 = (1'h0);
  reg [(2'h2):(1'h0)] reg843 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg842 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg840 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg836 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg835 = (1'h0);
  reg [(2'h2):(1'h0)] reg834 = (1'h0);
  reg [(5'h16):(1'h0)] forvar833 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg830 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg828 = (1'h0);
  assign y = {wire1312,
                 wire1167,
                 wire821,
                 wire823,
                 wire824,
                 wire825,
                 wire862,
                 wire994,
                 wire1169,
                 wire1170,
                 wire1171,
                 wire1190,
                 wire1191,
                 wire1288,
                 wire1290,
                 wire1292,
                 reg1311,
                 reg1310,
                 reg1308,
                 reg1307,
                 reg1304,
                 reg1303,
                 reg1300,
                 reg1299,
                 reg1296,
                 reg1187,
                 reg1186,
                 reg1185,
                 reg1179,
                 reg1183,
                 reg1177,
                 reg1175,
                 reg1174,
                 reg1172,
                 reg1020,
                 reg1019,
                 reg1017,
                 reg1014,
                 reg1011,
                 reg1010,
                 reg1008,
                 reg1007,
                 reg1005,
                 reg1003,
                 reg999,
                 reg998,
                 reg826,
                 reg827,
                 reg829,
                 reg831,
                 reg832,
                 reg837,
                 reg838,
                 reg839,
                 reg841,
                 reg846,
                 reg848,
                 reg851,
                 reg852,
                 reg854,
                 reg857,
                 reg858,
                 reg859,
                 reg861,
                 reg1309,
                 forvar1306,
                 reg1305,
                 forvar1302,
                 forvar1301,
                 reg1298,
                 reg1297,
                 forvar1295,
                 forvar1294,
                 reg1189,
                 reg1188,
                 reg1184,
                 reg1182,
                 reg1181,
                 reg1180,
                 forvar1179,
                 reg1178,
                 reg1176,
                 forvar1173,
                 reg1024,
                 reg1023,
                 reg1022,
                 reg1021,
                 reg1018,
                 reg1016,
                 reg1015,
                 reg1013,
                 reg1012,
                 reg1009,
                 reg1006,
                 reg1004,
                 reg1002,
                 reg1001,
                 forvar1000,
                 forvar997,
                 reg996,
                 reg860,
                 reg856,
                 reg855,
                 forvar853,
                 reg850,
                 reg849,
                 forvar847,
                 reg845,
                 reg844,
                 reg833,
                 forvar826,
                 reg843,
                 reg842,
                 reg840,
                 reg836,
                 reg835,
                 reg834,
                 forvar833,
                 reg830,
                 reg828,
                 (1'h0)};
  module709 #() modinst822 (.y(wire821), .wire713(wire708), .wire712(wire704), .clk(clk), .wire711(wire707), .wire710(wire705));
  assign wire823 = wire707[(1'h0):(1'h0)];
  assign wire824 = $signed(((^~(&wire821[(1'h1):(1'h1)])) <<< ($signed(wire823) ?
                       wire707[(2'h2):(1'h0)] : wire706)));
  assign wire825 = ((~&wire706) ?
                       (wire708 && wire705) : wire823[(3'h5):(1'h1)]);
  always
    @(posedge clk) begin
      if ((($unsigned(wire706[(4'h9):(2'h3)]) << (~{$signed(wire704)})) ^~ (|wire708)))
        begin
          if ($unsigned(((($unsigned(wire704) ^~ (wire823 == wire824)) ~^ wire706) ?
              $signed(((wire705 ? wire823 : wire708) | {wire707,
                  wire706})) : wire821)))
            begin
              reg826 <= wire825;
              reg827 <= wire704[(4'hc):(4'h9)];
              reg828 = wire821[(1'h0):(1'h0)];
              reg829 <= (wire823 ?
                  $unsigned(wire707[(4'ha):(4'h8)]) : (wire707[(4'he):(3'h7)] ?
                      ($unsigned({wire706,
                          wire708}) ^~ reg826[(1'h0):(1'h0)]) : ($signed((reg826 >> wire824)) ?
                          (8'hb9) : (((8'ha0) == wire707) ^ $unsigned(wire706)))));
              reg830 = wire708;
            end
          else
            begin
              reg828 = (((wire821[(1'h0):(1'h0)] != wire825) ?
                      reg827[(4'ha):(1'h0)] : $unsigned((((7'h4a) > reg826) && $unsigned(wire824)))) ?
                  ((^{(reg829 << reg826),
                      reg828}) & ((-wire825[(2'h3):(1'h0)]) ?
                      wire705 : {wire708[(4'ha):(3'h7)],
                          (~|wire821)})) : (|{reg828[(4'h8):(1'h0)]}));
              reg829 <= wire824[(2'h3):(2'h3)];
              reg831 <= $signed({(&({wire821, (8'ha3)} ? reg826 : wire823)),
                  (~|$unsigned(wire821[(1'h1):(1'h1)]))});
              reg832 <= reg826;
            end
          for (forvar833 = (1'h0); (forvar833 < (1'h0)); forvar833 = (forvar833 + (1'h1)))
            begin
              reg834 = (({$unsigned((^reg832)),
                          ((reg826 != reg826) ~^ (reg826 << wire705))} ?
                      (($signed((8'hb8)) | reg831) - (8'h9d)) : ($signed((reg832 ?
                              reg828 : (8'ha0))) ?
                          $signed((wire821 | forvar833)) : forvar833[(5'h13):(4'he)])) ?
                  ($unsigned(reg827) != $unsigned(reg826)) : wire706[(5'h11):(4'hb)]);
              reg835 = $unsigned(reg830);
              reg836 = $unsigned($signed({reg834}));
            end
          reg837 <= $signed(wire824[(3'h4):(2'h3)]);
          if ($unsigned($signed($unsigned($signed((8'hb8))))))
            begin
              reg838 <= $signed(reg829[(2'h3):(1'h0)]);
              reg839 <= (8'hb6);
              reg840 = wire708[(4'hc):(1'h0)];
              reg841 <= (-(^~((+(reg828 == reg838)) ?
                  $signed((reg835 != reg832)) : reg828[(4'ha):(4'h9)])));
            end
          else
            begin
              reg838 <= (wire704[(3'h7):(3'h6)] ?
                  (reg841 | {(reg840[(2'h3):(1'h1)] & $unsigned((8'hb2))),
                      {(-reg828), wire707}}) : ({$unsigned((wire707 ?
                          reg839 : wire824))} - ((reg829 > wire823[(2'h2):(1'h1)]) ?
                      (((8'ha2) >= reg834) ?
                          (wire706 >>> forvar833) : (wire823 ?
                              reg828 : wire825)) : reg838)));
              reg839 <= $signed((8'ha8));
              reg840 = {(!{($signed(reg831) ?
                          $unsigned(reg835) : (reg838 == reg839))}),
                  (~$signed({forvar833}))};
              reg841 <= $unsigned(wire708[(3'h7):(3'h6)]);
              reg842 = wire707[(2'h2):(1'h0)];
            end
          reg843 = (^~(|$signed(((reg831 ?
              reg834 : forvar833) <= reg826[(3'h4):(1'h0)]))));
        end
      else
        begin
          for (forvar826 = (1'h0); (forvar826 < (2'h3)); forvar826 = (forvar826 + (1'h1)))
            begin
              reg828 = (-reg828[(4'hb):(3'h6)]);
              reg830 = (wire705 ? reg836 : $unsigned(reg842));
              reg831 <= reg829;
            end
          if ((($signed(($unsigned(reg841) || $unsigned(reg835))) ?
              (reg834 ?
                  ((8'ha5) ?
                      wire708[(4'hb):(3'h7)] : reg832[(4'hf):(4'ha)]) : $unsigned(wire704)) : (!(reg827[(4'h8):(1'h1)] <<< reg832[(4'ha):(3'h6)]))) && $signed($signed(reg838[(4'hd):(3'h7)]))))
            begin
              reg833 = (($unsigned($unsigned((reg836 < (7'h43)))) - $unsigned(((~^(8'ha8)) - (&reg837)))) || {reg828[(3'h7):(1'h1)]});
              reg837 <= reg836[(4'ha):(3'h6)];
              reg840 = (!wire708);
            end
          else
            begin
              reg832 <= (8'hae);
              reg837 <= ($signed(wire707[(5'h11):(1'h0)]) ?
                  (reg835[(3'h6):(3'h4)] ?
                      wire821[(1'h1):(1'h1)] : (forvar833[(1'h1):(1'h1)] >>> $signed(reg835))) : (~wire707[(2'h3):(1'h1)]));
              reg840 = $unsigned({((~^$signed((7'h43))) - $signed((reg842 && reg832))),
                  (^~($signed(wire706) >>> {reg830}))});
              reg842 = ((({(reg828 && wire706),
                      (+reg832)} * $unsigned(reg828)) ^ (!(&(wire705 ~^ forvar826)))) ?
                  wire704[(4'hc):(2'h2)] : {wire825,
                      ($signed($unsigned(wire705)) != $unsigned((~|reg826)))});
              reg843 = wire704[(2'h3):(2'h3)];
            end
          reg844 = $unsigned(($unsigned(($signed((8'hb7)) + (reg827 >= wire821))) ?
              (~{{reg842, reg838}, (8'hbc)}) : $signed(reg842)));
        end
    end
  always
    @(posedge clk) begin
      reg845 = (-reg841[(3'h7):(3'h6)]);
      reg846 <= (^wire821[(2'h2):(1'h1)]);
      for (forvar847 = (1'h0); (forvar847 < (1'h1)); forvar847 = (forvar847 + (1'h1)))
        begin
          reg848 <= $signed(reg837);
          reg849 = ((8'hba) ? wire707[(4'ha):(4'h8)] : wire704);
          if (($signed(reg829) || (wire705 && ($signed($signed(reg827)) ?
              ((~&wire707) != ((7'h4a) ? reg832 : (8'hb8))) : reg826))))
            begin
              reg850 = $signed((!$signed(reg849[(1'h0):(1'h0)])));
            end
          else
            begin
              reg851 <= (^$unsigned($signed((reg848 < (|reg841)))));
              reg852 <= $unsigned((~$signed({((8'ha0) * reg849)})));
            end
          for (forvar853 = (1'h0); (forvar853 < (1'h0)); forvar853 = (forvar853 + (1'h1)))
            begin
              reg854 <= {{reg829[(2'h3):(1'h1)],
                      $unsigned($signed((wire825 ? forvar853 : reg848)))},
                  ($signed((!(reg852 & reg826))) - ($signed($signed(wire704)) ?
                      $signed({reg850, reg848}) : (wire821 ?
                          ((8'h9c) + (8'hb4)) : wire821)))};
              reg855 = wire708[(3'h6):(3'h6)];
            end
          if ((reg826[(2'h3):(2'h3)] ?
              wire706[(5'h15):(2'h3)] : (reg831 ?
                  (wire704[(3'h4):(2'h3)] ?
                      reg831[(5'h17):(1'h0)] : $signed(reg855[(4'h9):(2'h2)])) : $signed($signed(wire704[(3'h4):(2'h3)])))))
            begin
              reg856 = {wire705, $signed((8'hb4))};
              reg857 <= wire708;
              reg858 <= ((((((7'h47) ?
                          reg855 : reg850) ^ $unsigned(wire821)) << {(reg829 ?
                              reg848 : reg852)}) ?
                      $unsigned(wire705[(3'h5):(3'h5)]) : $signed(reg855)) ?
                  (+(+$signed((wire825 + reg846)))) : wire704[(3'h5):(2'h2)]);
              reg859 <= reg854[(1'h1):(1'h0)];
            end
          else
            begin
              reg856 = $signed(($unsigned(wire823) ?
                  $signed($unsigned(reg831[(4'h9):(3'h7)])) : reg855[(4'h9):(1'h0)]));
              reg857 <= {reg854,
                  $signed((($unsigned(reg838) ?
                      reg858 : $unsigned((8'hb1))) - reg846))};
              reg858 <= {wire821[(1'h0):(1'h0)]};
              reg860 = $signed(($unsigned(reg850[(2'h2):(1'h0)]) ?
                  wire708 : reg839[(3'h4):(2'h3)]));
              reg861 <= $unsigned(reg839[(3'h7):(2'h3)]);
            end
        end
    end
  assign wire862 = $signed($signed((((~|wire821) ?
                           (7'h40) : (reg861 & wire708)) ?
                       reg838 : (~|wire825))));
  module863 #() modinst995 (.wire865(wire705), .wire867(reg837), .wire864(reg852), .y(wire994), .clk(clk), .wire866(reg832));
  always
    @(posedge clk) begin
      reg996 = reg827;
      for (forvar997 = (1'h0); (forvar997 < (2'h3)); forvar997 = (forvar997 + (1'h1)))
        begin
          reg998 <= (reg838 ?
              $signed($signed(reg858)) : {$signed((reg841[(2'h2):(2'h2)] ?
                      (^~wire823) : (wire994 < (8'h9d)))),
                  reg839[(4'hb):(2'h3)]});
        end
      reg999 <= {reg858[(4'h9):(4'h9)],
          (({$signed(wire823), $unsigned((8'hac))} ?
                  $signed($unsigned((8'hb6))) : (+(reg996 >= wire821))) ?
              reg851[(2'h3):(1'h0)] : wire707[(4'ha):(4'h9)])};
      for (forvar1000 = (1'h0); (forvar1000 < (2'h3)); forvar1000 = (forvar1000 + (1'h1)))
        begin
          reg1001 = (((~^(8'hb2)) >>> $unsigned({reg827[(4'hd):(4'h8)]})) ?
              $signed(wire824[(3'h7):(3'h7)]) : wire706);
          reg1002 = reg852;
        end
    end
  always
    @(posedge clk) begin
      if ((8'h9f))
        begin
          if ($signed($signed($signed($unsigned((wire821 <<< wire705))))))
            begin
              reg1003 <= {((7'h49) != $signed(reg852)),
                  ($unsigned(reg831[(5'h12):(5'h10)]) || (((&reg846) ?
                      wire706[(1'h0):(1'h0)] : wire705[(5'h16):(3'h4)]) - (7'h41)))};
              reg1004 = reg859[(3'h5):(2'h3)];
              reg1005 <= reg852[(1'h0):(1'h0)];
              reg1006 = (7'h49);
              reg1007 <= (reg826 ?
                  {{{(wire706 && (8'haf))}, (^(reg857 ^~ reg858))},
                      reg838[(3'h5):(3'h4)]} : $signed(wire821[(2'h2):(1'h0)]));
            end
          else
            begin
              reg1003 <= reg1006;
              reg1005 <= wire824[(3'h5):(1'h1)];
              reg1007 <= reg841[(2'h2):(1'h0)];
              reg1008 <= ((reg839 || ($signed((reg1006 | wire825)) ~^ $unsigned(reg1003[(4'h8):(2'h3)]))) ?
                  (reg1003 <<< $signed((wire825[(2'h2):(1'h0)] ?
                      reg861[(2'h2):(1'h1)] : wire705))) : reg999[(4'ha):(2'h3)]);
              reg1009 = $unsigned($signed(reg841));
            end
          if (reg857)
            begin
              reg1010 <= $unsigned(({(|((8'ha1) ? wire706 : reg839))} ?
                  (+reg857[(1'h1):(1'h1)]) : (~|(!reg829))));
              reg1011 <= ($signed(reg859[(1'h1):(1'h0)]) ?
                  reg827[(1'h0):(1'h0)] : wire704);
              reg1012 = $unsigned(reg1008);
              reg1013 = wire708[(2'h3):(1'h1)];
            end
          else
            begin
              reg1012 = ($unsigned({reg1011}) ?
                  $unsigned(reg831) : {($signed($signed(reg829)) ?
                          (^(reg1006 >= (8'haf))) : ((^reg1005) ?
                              $signed(wire708) : (reg1007 ? reg852 : reg1003))),
                      {{((8'hba) ? reg1008 : reg1012)}}});
              reg1014 <= reg861[(2'h3):(1'h0)];
              reg1015 = ((~^({reg826,
                  (reg1005 && reg827)} + wire823[(1'h1):(1'h0)])) & ({reg857[(4'h8):(2'h3)],
                      ($unsigned(reg1006) ? reg838[(1'h0):(1'h0)] : (8'hb7))} ?
                  $signed(reg829) : $signed(($signed(wire708) ^~ (~^(8'hae))))));
              reg1016 = reg851;
            end
          if ((~reg1004))
            begin
              reg1017 <= reg826;
            end
          else
            begin
              reg1018 = $unsigned($signed((wire862[(1'h1):(1'h1)] ?
                  (wire994 && (!wire708)) : {reg852[(4'he):(4'h9)],
                      (reg1013 <= reg1006)})));
              reg1019 <= {wire823[(4'hd):(4'hb)]};
            end
          reg1020 <= $unsigned($signed($signed((reg831 >= (reg857 ?
              reg1009 : reg1009)))));
          reg1021 = $signed((reg1012[(2'h2):(1'h1)] * (reg1004 ?
              {((8'hb2) <<< reg857)} : $signed($signed(reg1009)))));
        end
      else
        begin
          reg1003 <= $signed($unsigned($unsigned($unsigned($unsigned(reg1017)))));
          if ((!((((8'hae) ~^ (&wire862)) ?
              (!$signed((8'ha5))) : $unsigned((wire704 ?
                  reg831 : reg1013))) << (((~reg829) ?
              $signed(wire823) : reg1005) | ($unsigned((8'hb2)) | {reg1007,
              reg1017})))))
            begin
              reg1004 = (reg1018[(5'h13):(3'h4)] <<< reg827);
              reg1005 <= $signed(($unsigned((^~{reg837, reg854})) ?
                  reg861 : $unsigned($unsigned($signed((8'haf))))));
              reg1007 <= (reg826 ?
                  $unsigned(reg848) : (+(reg1017[(5'h17):(3'h6)] ?
                      $unsigned((wire824 | reg854)) : (+wire994))));
              reg1009 = ((reg1015 < $unsigned({$signed(reg859)})) | $signed((~^$signed(reg1004[(1'h1):(1'h1)]))));
              reg1010 <= wire994;
            end
          else
            begin
              reg1005 <= reg1014[(3'h5):(2'h3)];
              reg1006 = $unsigned($signed((8'hb8)));
              reg1009 = $unsigned($unsigned($signed($signed(reg999))));
              reg1010 <= $unsigned(((&wire707) << (~$signed((^~reg1007)))));
              reg1011 <= (-reg1007);
            end
          if (reg829[(4'hc):(3'h7)])
            begin
              reg1014 <= $signed(reg826[(3'h4):(3'h4)]);
              reg1017 <= $unsigned((($signed({reg1006}) ?
                  ((^~(7'h48)) >> wire821) : {$unsigned(reg1011),
                      $unsigned(reg1012)}) <<< (~^(~&{(8'hbc), reg831}))));
              reg1018 = (8'hbf);
              reg1021 = reg1009;
              reg1022 = reg829;
            end
          else
            begin
              reg1014 <= {(8'ha2)};
              reg1015 = (!reg859[(2'h3):(2'h2)]);
              reg1017 <= $unsigned(wire706);
              reg1019 <= reg852[(3'h4):(2'h2)];
            end
        end
      reg1023 = (!(~^reg1020));
      reg1024 = (!(-$unsigned($signed((reg826 ? wire825 : reg1020)))));
    end
  module1025 #() modinst1168 (.wire1030(reg846), .clk(clk), .wire1026(reg841), .wire1028(wire862), .wire1027(reg838), .y(wire1167), .wire1029(reg857));
  assign wire1169 = wire823;
  assign wire1170 = $signed(wire824);
  assign wire1171 = (+(~(~|(7'h49))));
  always
    @(posedge clk) begin
      reg1172 <= wire705[(3'h7):(3'h4)];
      for (forvar1173 = (1'h0); (forvar1173 < (2'h2)); forvar1173 = (forvar1173 + (1'h1)))
        begin
          reg1174 <= (((^({wire704} != {reg852, reg1005})) ?
                  wire1170[(2'h2):(2'h2)] : {{(~|reg848), $signed((8'hbb))}}) ?
              $signed({((wire707 ? (8'hbc) : (7'h48)) << (reg841 ?
                      reg854 : wire707))}) : $signed(($unsigned($signed(wire825)) << ((8'ha7) - $unsigned(reg832)))));
          reg1175 <= wire862;
          reg1176 = $signed($signed((^reg1175)));
          reg1177 <= (({(^reg1007),
              $signed(reg1017)} << $signed($unsigned($signed(reg861)))) << {reg854});
        end
      if ($signed($unsigned(reg1172[(2'h3):(1'h0)])))
        begin
          reg1178 = $signed((~|(-($signed(wire824) ?
              (wire705 ? wire824 : (8'h9c)) : reg1005[(5'h12):(4'ha)]))));
          for (forvar1179 = (1'h0); (forvar1179 < (2'h3)); forvar1179 = (forvar1179 + (1'h1)))
            begin
              reg1180 = (reg826 ? wire994 : (^$signed({reg1178})));
              reg1181 = wire823[(2'h3):(2'h2)];
              reg1182 = ($unsigned((~|$signed({reg1172}))) <<< (-$signed((~^$unsigned((8'hbc))))));
              reg1183 <= $signed($unsigned(reg1175));
              reg1184 = (($signed($unsigned((|forvar1179))) ?
                  $signed(($unsigned(reg1174) > (reg1017 >= wire704))) : ((reg1020 ?
                          (~^reg1010) : $signed(reg999)) ?
                      reg1182[(3'h4):(1'h0)] : $unsigned((~|wire994)))) >= ({((reg1008 ?
                              (8'ha6) : wire1170) ?
                          $signed(reg852) : $signed((8'hb7)))} ?
                  (((reg1174 ? reg827 : reg861) ?
                          $unsigned(reg826) : $signed((8'h9f))) ?
                      $signed((~|reg1014)) : ($signed(reg1181) ?
                          (reg1008 ?
                              wire706 : reg858) : (reg861 | reg1017))) : (|$signed({reg1007,
                      reg846}))));
            end
        end
      else
        begin
          reg1179 <= (wire823 > {$unsigned($signed((reg1177 ?
                  reg829 : reg1017))),
              (($signed(reg998) ?
                      reg998[(4'hc):(4'h8)] : (reg841 ? reg1017 : reg848)) ?
                  reg831[(4'hf):(3'h4)] : reg857[(2'h2):(1'h0)])});
          if (reg1182[(4'ha):(1'h1)])
            begin
              reg1183 <= wire821[(1'h1):(1'h1)];
              reg1185 <= $unsigned(($signed($signed(reg839[(4'he):(1'h0)])) + (-{(|reg1020),
                  (~&forvar1173)})));
              reg1186 <= $signed(reg846);
              reg1187 <= reg838;
              reg1188 = $unsigned((reg859 > {$unsigned($unsigned(reg1011)),
                  $unsigned((-forvar1173))}));
            end
          else
            begin
              reg1183 <= $unsigned($signed((7'h49)));
              reg1185 <= reg1179;
            end
        end
    end
  always
    @(posedge clk) begin
      reg1189 = (!(+{((!reg827) ?
              $unsigned(reg1175) : reg839[(4'hd):(4'h9)])}));
    end
  assign wire1190 = (reg829[(4'h8):(1'h0)] ?
                        (8'ha2) : $unsigned((-(~|wire862[(3'h4):(1'h0)]))));
  assign wire1191 = (~(7'h42));
  module1192 #() modinst1289 (.wire1195(reg839), .clk(clk), .wire1193(reg857), .wire1196(reg1014), .y(wire1288), .wire1197(reg831), .wire1194(reg848));
  module863 #() modinst1291 (.clk(clk), .wire866(reg1003), .wire867(reg829), .wire864(reg1185), .wire865(reg1011), .y(wire1290));
  module709 #() modinst1293 (.wire712(reg827), .y(wire1292), .wire710(reg858), .wire711(reg859), .clk(clk), .wire713(wire994));
  always
    @(posedge clk) begin
      for (forvar1294 = (1'h0); (forvar1294 < (1'h0)); forvar1294 = (forvar1294 + (1'h1)))
        begin
          for (forvar1295 = (1'h0); (forvar1295 < (1'h0)); forvar1295 = (forvar1295 + (1'h1)))
            begin
              reg1296 <= ($unsigned(reg1014[(5'h13):(4'h9)]) <= (reg839[(4'hd):(3'h7)] ?
                  (8'ha3) : $signed(reg829[(4'hc):(3'h6)])));
              reg1297 = (wire705 ?
                  $unsigned((+$signed((reg838 >= reg1179)))) : (($signed(((8'hb2) ?
                          reg1010 : (8'hb5))) ?
                      $signed(reg1179[(2'h3):(2'h2)]) : {reg1005}) <<< (^~wire704)));
              reg1298 = reg1010[(4'ha):(1'h1)];
            end
        end
      reg1299 <= ((~|$signed((wire1288[(2'h2):(2'h2)] + {reg998,
          reg827}))) ~^ ($signed((^$unsigned(reg1007))) | $signed(((reg846 | reg1020) < $signed(reg1179)))));
      reg1300 <= (reg858[(4'hb):(4'h8)] ?
          ((reg1007 ? (~reg846) : $unsigned(((8'hb9) ? reg1175 : wire1171))) ?
              (8'hb0) : (((reg848 ? reg1014 : wire862) ?
                      (+reg861) : (reg1010 ? reg846 : reg1020)) ?
                  reg1010[(3'h5):(1'h0)] : {(wire994 ?
                          reg858 : reg1187)})) : (~$unsigned((8'hb7))));
      for (forvar1301 = (1'h0); (forvar1301 < (1'h0)); forvar1301 = (forvar1301 + (1'h1)))
        begin
          for (forvar1302 = (1'h0); (forvar1302 < (2'h3)); forvar1302 = (forvar1302 + (1'h1)))
            begin
              reg1303 <= reg1179[(2'h3):(1'h1)];
              reg1304 <= reg1175;
              reg1305 = (7'h47);
            end
          for (forvar1306 = (1'h0); (forvar1306 < (1'h1)); forvar1306 = (forvar1306 + (1'h1)))
            begin
              reg1307 <= wire706[(5'h10):(4'hc)];
              reg1308 <= (reg1183[(4'h9):(3'h7)] - $signed($signed($unsigned({(8'hb8),
                  wire707}))));
              reg1309 = reg1008;
              reg1310 <= $signed(reg831);
            end
          reg1311 <= ({(~((8'hbc) <<< (8'hb6)))} ?
              ($signed($unsigned(reg826)) ?
                  (~((forvar1306 ?
                      (8'h9f) : reg1179) + (forvar1306 | reg1308))) : ($signed((reg1298 ?
                          reg838 : wire862)) ?
                      $unsigned((~&reg839)) : $unsigned((reg832 ?
                          (8'haa) : reg841)))) : reg1185[(4'hb):(1'h0)]);
        end
    end
  assign wire1312 = (^reg1175);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module279
#(parameter param649 = (((8'hb2) ? ((((8'h9e) ? (8'ha6) : (8'hb8)) ? ((8'hb5) >>> (8'ha0)) : (+(8'hb0))) && (^~(|(7'h40)))) : {(-{(8'hb0), (8'hac)})}) ? {((~((7'h48) && (8'hac))) | (((8'hb2) ? (8'ha3) : (8'had)) == (~(8'ha3)))), (~|{((8'hac) >> (7'h47))})} : (((((8'ha3) ? (8'hb3) : (8'hba)) ? (~|(8'hb9)) : ((8'hb7) ? (8'h9e) : (8'ha3))) ? {(8'h9e)} : {((8'hb3) != (7'h49))}) <= (({(8'hb9), (8'ha4)} ? {(8'h9f)} : ((8'hbc) <= (7'h41))) - (((8'haf) ? (7'h49) : (8'hb9)) << (^~(8'ha3)))))))
(y, clk, wire280, wire281, wire282, wire283, wire284);
  output wire [(32'h766):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire280;
  input wire [(4'he):(1'h0)] wire281;
  input wire signed [(4'hb):(1'h0)] wire282;
  input wire [(5'h16):(1'h0)] wire283;
  input wire signed [(5'h11):(1'h0)] wire284;
  wire signed [(4'ha):(1'h0)] wire630;
  wire [(4'he):(1'h0)] wire624;
  wire signed [(5'h18):(1'h0)] wire622;
  wire [(5'h16):(1'h0)] wire306;
  wire signed [(4'hd):(1'h0)] wire307;
  wire [(4'he):(1'h0)] wire341;
  wire signed [(4'hf):(1'h0)] wire348;
  wire signed [(4'hf):(1'h0)] wire392;
  wire signed [(4'hb):(1'h0)] wire393;
  wire signed [(3'h4):(1'h0)] wire426;
  reg signed [(4'h8):(1'h0)] reg646 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg645 = (1'h0);
  reg [(5'h18):(1'h0)] reg642 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg641 = (1'h0);
  reg [(3'h6):(1'h0)] reg638 = (1'h0);
  reg [(4'he):(1'h0)] reg637 = (1'h0);
  reg [(4'he):(1'h0)] reg634 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg632 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg631 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg629 = (1'h0);
  reg [(2'h2):(1'h0)] reg388 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg387 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg386 = (1'h0);
  reg [(5'h16):(1'h0)] reg385 = (1'h0);
  reg [(4'h8):(1'h0)] reg376 = (1'h0);
  reg [(5'h10):(1'h0)] reg381 = (1'h0);
  reg [(2'h3):(1'h0)] reg378 = (1'h0);
  reg [(4'hf):(1'h0)] reg373 = (1'h0);
  reg [(3'h5):(1'h0)] reg370 = (1'h0);
  reg [(5'h14):(1'h0)] reg369 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg368 = (1'h0);
  reg [(2'h3):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg352 = (1'h0);
  reg [(4'hb):(1'h0)] reg363 = (1'h0);
  reg [(5'h14):(1'h0)] reg362 = (1'h0);
  reg [(5'h16):(1'h0)] reg361 = (1'h0);
  reg [(4'hf):(1'h0)] reg360 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg356 = (1'h0);
  reg [(4'hb):(1'h0)] reg355 = (1'h0);
  reg [(5'h18):(1'h0)] reg349 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg347 = (1'h0);
  reg [(4'ha):(1'h0)] reg343 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg342 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg340 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg337 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg335 = (1'h0);
  reg [(3'h4):(1'h0)] reg331 = (1'h0);
  reg [(3'h7):(1'h0)] reg329 = (1'h0);
  reg [(2'h3):(1'h0)] reg327 = (1'h0);
  reg [(3'h7):(1'h0)] reg326 = (1'h0);
  reg [(5'h13):(1'h0)] reg322 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg321 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg319 = (1'h0);
  reg [(5'h13):(1'h0)] reg315 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg314 = (1'h0);
  reg [(5'h10):(1'h0)] reg309 = (1'h0);
  reg [(4'h9):(1'h0)] reg305 = (1'h0);
  reg [(5'h15):(1'h0)] reg302 = (1'h0);
  reg [(5'h10):(1'h0)] reg301 = (1'h0);
  reg [(4'hf):(1'h0)] reg299 = (1'h0);
  reg [(5'h10):(1'h0)] reg294 = (1'h0);
  reg [(5'h13):(1'h0)] reg291 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg290 = (1'h0);
  reg [(3'h7):(1'h0)] reg289 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg288 = (1'h0);
  reg [(4'hc):(1'h0)] reg287 = (1'h0);
  reg [(5'h12):(1'h0)] reg648 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg647 = (1'h0);
  reg [(5'h17):(1'h0)] reg644 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar643 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar640 = (1'h0);
  reg [(4'he):(1'h0)] reg639 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg636 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar635 = (1'h0);
  reg [(5'h13):(1'h0)] forvar633 = (1'h0);
  reg [(2'h3):(1'h0)] reg628 = (1'h0);
  reg [(5'h11):(1'h0)] forvar627 = (1'h0);
  reg [(3'h7):(1'h0)] reg626 = (1'h0);
  reg [(5'h12):(1'h0)] reg625 = (1'h0);
  reg [(5'h13):(1'h0)] reg391 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg390 = (1'h0);
  reg signed [(4'he):(1'h0)] reg389 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar384 = (1'h0);
  reg [(5'h10):(1'h0)] reg383 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar382 = (1'h0);
  reg [(5'h12):(1'h0)] reg380 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg379 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg377 = (1'h0);
  reg [(5'h18):(1'h0)] forvar376 = (1'h0);
  reg [(3'h6):(1'h0)] reg375 = (1'h0);
  reg [(4'ha):(1'h0)] reg374 = (1'h0);
  reg [(5'h14):(1'h0)] reg372 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg367 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg366 = (1'h0);
  reg [(5'h14):(1'h0)] reg365 = (1'h0);
  reg [(5'h18):(1'h0)] forvar361 = (1'h0);
  reg [(4'he):(1'h0)] reg357 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar349 = (1'h0);
  reg signed [(4'he):(1'h0)] reg359 = (1'h0);
  reg [(4'he):(1'h0)] reg358 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar357 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg354 = (1'h0);
  reg [(4'h9):(1'h0)] reg353 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar352 = (1'h0);
  reg [(5'h11):(1'h0)] reg351 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg350 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg346 = (1'h0);
  reg [(4'h8):(1'h0)] reg345 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar344 = (1'h0);
  reg [(3'h6):(1'h0)] forvar335 = (1'h0);
  reg [(5'h17):(1'h0)] reg339 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg338 = (1'h0);
  reg [(5'h10):(1'h0)] reg336 = (1'h0);
  reg [(5'h17):(1'h0)] reg334 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg333 = (1'h0);
  reg [(4'ha):(1'h0)] reg332 = (1'h0);
  reg [(4'hc):(1'h0)] reg330 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar328 = (1'h0);
  reg [(5'h12):(1'h0)] reg325 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar324 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg320 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg318 = (1'h0);
  reg [(3'h5):(1'h0)] forvar317 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar316 = (1'h0);
  reg [(4'hf):(1'h0)] reg313 = (1'h0);
  reg [(2'h3):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg311 = (1'h0);
  reg [(3'h7):(1'h0)] forvar310 = (1'h0);
  reg [(3'h6):(1'h0)] reg308 = (1'h0);
  reg [(4'hf):(1'h0)] reg304 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg303 = (1'h0);
  reg [(3'h5):(1'h0)] forvar300 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg298 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg297 = (1'h0);
  reg [(3'h7):(1'h0)] reg296 = (1'h0);
  reg [(4'h8):(1'h0)] forvar295 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg293 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg292 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar286 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar285 = (1'h0);
  assign y = {wire630,
                 wire624,
                 wire622,
                 wire306,
                 wire307,
                 wire341,
                 wire348,
                 wire392,
                 wire393,
                 wire426,
                 reg646,
                 reg645,
                 reg642,
                 reg641,
                 reg638,
                 reg637,
                 reg634,
                 reg632,
                 reg631,
                 reg629,
                 reg388,
                 reg387,
                 reg386,
                 reg385,
                 reg376,
                 reg381,
                 reg378,
                 reg373,
                 reg370,
                 reg369,
                 reg368,
                 reg364,
                 reg352,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 reg356,
                 reg355,
                 reg349,
                 reg347,
                 reg343,
                 reg342,
                 reg340,
                 reg337,
                 reg335,
                 reg331,
                 reg329,
                 reg327,
                 reg326,
                 reg322,
                 reg321,
                 reg319,
                 reg315,
                 reg314,
                 reg309,
                 reg305,
                 reg302,
                 reg301,
                 reg299,
                 reg294,
                 reg291,
                 reg290,
                 reg289,
                 reg288,
                 reg287,
                 reg648,
                 reg647,
                 reg644,
                 forvar643,
                 forvar640,
                 reg639,
                 reg636,
                 forvar635,
                 forvar633,
                 reg628,
                 forvar627,
                 reg626,
                 reg625,
                 reg391,
                 reg390,
                 reg389,
                 forvar384,
                 reg383,
                 forvar382,
                 reg380,
                 reg379,
                 reg377,
                 forvar376,
                 reg375,
                 reg374,
                 reg372,
                 reg371,
                 reg367,
                 reg366,
                 reg365,
                 forvar361,
                 reg357,
                 forvar349,
                 reg359,
                 reg358,
                 forvar357,
                 reg354,
                 reg353,
                 forvar352,
                 reg351,
                 reg350,
                 reg346,
                 reg345,
                 forvar344,
                 forvar335,
                 reg339,
                 reg338,
                 reg336,
                 reg334,
                 reg333,
                 reg332,
                 reg330,
                 forvar328,
                 reg325,
                 forvar324,
                 reg323,
                 reg320,
                 reg318,
                 forvar317,
                 forvar316,
                 reg313,
                 reg312,
                 reg311,
                 forvar310,
                 reg308,
                 reg304,
                 reg303,
                 forvar300,
                 reg298,
                 reg297,
                 reg296,
                 forvar295,
                 reg293,
                 reg292,
                 forvar286,
                 forvar285,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar285 = (1'h0); (forvar285 < (2'h3)); forvar285 = (forvar285 + (1'h1)))
        begin
          for (forvar286 = (1'h0); (forvar286 < (2'h3)); forvar286 = (forvar286 + (1'h1)))
            begin
              reg287 <= (^wire282);
              reg288 <= (($signed(((wire284 || forvar285) ?
                      (^wire283) : (~wire283))) <<< {forvar285[(3'h5):(2'h2)],
                      $signed((8'ha5))}) ?
                  reg287 : $unsigned((^~(~&$signed(reg287)))));
              reg289 <= reg288[(3'h5):(3'h5)];
              reg290 <= $unsigned($signed(wire280));
            end
          if (($unsigned($unsigned(((wire281 <= reg288) ?
                  (|wire281) : forvar286))) ?
              wire284[(5'h10):(4'hb)] : (!{$unsigned((~^wire283))})))
            begin
              reg291 <= (!$unsigned(reg289));
              reg292 = {$unsigned($signed($unsigned((forvar285 ?
                      (7'h47) : reg288))))};
            end
          else
            begin
              reg292 = {(~(reg289[(2'h2):(1'h1)] ?
                      wire283[(4'hb):(3'h5)] : wire284)),
                  $signed((-(~(~wire281))))};
              reg293 = {reg291};
            end
          reg294 <= $signed(wire284);
          for (forvar295 = (1'h0); (forvar295 < (1'h0)); forvar295 = (forvar295 + (1'h1)))
            begin
              reg296 = {forvar285[(1'h1):(1'h0)], wire282[(3'h6):(3'h4)]};
              reg297 = forvar285;
              reg298 = $unsigned((reg290[(3'h4):(2'h3)] ?
                  ($signed((reg296 ?
                      wire282 : (7'h40))) || ($signed(forvar285) >>> reg290)) : {{{reg292}}}));
              reg299 <= (~&(($unsigned(wire281[(4'h8):(2'h3)]) ?
                      {forvar285[(3'h4):(1'h1)], forvar286} : wire280) ?
                  (^~reg289) : (($unsigned(reg287) ?
                          (wire284 ?
                              forvar286 : reg298) : (reg293 << (8'hbb))) ?
                      $signed(((8'hb3) && forvar285)) : ((reg292 ?
                          reg292 : reg287) || (~|reg287)))));
            end
        end
      if ((~($signed(forvar295[(3'h7):(3'h6)]) ?
          (($unsigned(reg294) ?
                  reg290[(3'h6):(3'h4)] : (wire283 ? reg290 : reg287)) ?
              (~&$signed((8'ha1))) : ((reg293 ^ forvar286) ?
                  reg287[(1'h1):(1'h1)] : {forvar285})) : $signed($unsigned(reg287[(1'h1):(1'h1)])))))
        begin
          for (forvar300 = (1'h0); (forvar300 < (1'h0)); forvar300 = (forvar300 + (1'h1)))
            begin
              reg301 <= reg298;
            end
          reg302 <= reg289[(2'h3):(2'h3)];
          reg303 = {((reg287[(2'h2):(2'h2)] * (wire284[(1'h0):(1'h0)] ?
                      (wire281 - reg294) : (forvar286 ? (8'hba) : reg294))) ?
                  $signed(wire282[(1'h1):(1'h0)]) : forvar295[(2'h2):(2'h2)]),
              (forvar286 ? wire280[(4'h9):(2'h3)] : reg290[(3'h5):(1'h1)])};
          reg304 = $signed(reg299[(3'h4):(1'h0)]);
        end
      else
        begin
          for (forvar300 = (1'h0); (forvar300 < (2'h2)); forvar300 = (forvar300 + (1'h1)))
            begin
              reg303 = $unsigned(((^(~&$signed(wire284))) ?
                  $unsigned(reg303) : {$signed(reg301),
                      (~|((7'h43) == reg293))}));
              reg304 = (~&$unsigned((reg301[(3'h5):(3'h5)] <= forvar300)));
            end
          reg305 <= $signed((-($signed(forvar286) ^ (reg291[(4'hb):(3'h5)] <= reg288[(5'h12):(2'h3)]))));
        end
    end
  assign wire306 = $signed(($signed(reg299) ?
                       ($unsigned($signed(reg302)) ?
                           $unsigned({wire283}) : (&$signed((7'h48)))) : ((|reg287) ?
                           reg288[(2'h2):(2'h2)] : wire282[(1'h0):(1'h0)])));
  assign wire307 = ({$unsigned(reg294),
                       (7'h43)} == (((^(reg290 > wire281)) == wire283) ?
                       $unsigned(($unsigned(wire283) ?
                           (8'hb3) : (reg290 ?
                               reg299 : reg288))) : wire280[(1'h0):(1'h0)]));
  always
    @(posedge clk) begin
      if ($signed((reg299 >> wire280[(3'h4):(1'h1)])))
        begin
          reg308 = ({$signed(reg289[(1'h0):(1'h0)]),
              ((wire281 < (^~(8'hb9))) ?
                  wire280[(3'h7):(1'h0)] : reg302[(3'h7):(3'h5)])} > $signed(((^(wire280 ?
                  wire280 : reg305)) ?
              (~&(reg291 | wire280)) : wire307)));
        end
      else
        begin
          reg308 = reg291[(5'h13):(5'h11)];
          reg309 <= $unsigned((-{$unsigned((reg291 ? (7'h46) : (8'h9f)))}));
          for (forvar310 = (1'h0); (forvar310 < (3'h4)); forvar310 = (forvar310 + (1'h1)))
            begin
              reg311 = $unsigned($signed((~&$unsigned(wire307))));
              reg312 = {($signed($signed((wire280 >>> (8'ha9)))) ^~ $signed(reg309[(4'hf):(4'hf)])),
                  reg294[(2'h3):(1'h1)]};
              reg313 = {{((^$signed((8'hb6))) ?
                          reg302[(5'h11):(4'hc)] : (reg289 ?
                              (8'hae) : (~wire306))),
                      (wire306[(3'h5):(2'h3)] ?
                          wire281[(4'h8):(3'h5)] : reg302[(1'h1):(1'h1)])},
                  (((&(7'h47)) <<< (+reg305)) ?
                      {$signed({reg302, reg294})} : $signed(reg287))};
              reg314 <= (reg301 < reg302[(5'h13):(3'h4)]);
            end
          reg315 <= $signed($signed(wire283[(3'h5):(3'h5)]));
        end
      for (forvar316 = (1'h0); (forvar316 < (2'h2)); forvar316 = (forvar316 + (1'h1)))
        begin
          for (forvar317 = (1'h0); (forvar317 < (2'h3)); forvar317 = (forvar317 + (1'h1)))
            begin
              reg318 = (~reg287[(4'hb):(4'h8)]);
              reg319 <= $signed(wire284);
              reg320 = $signed($unsigned($signed(($unsigned(wire280) ?
                  reg305[(3'h5):(3'h5)] : $unsigned(reg319)))));
              reg321 <= (8'haa);
            end
          if (reg289[(3'h7):(1'h0)])
            begin
              reg322 <= $unsigned(reg299[(4'h9):(1'h0)]);
              reg323 = ((+(~$unsigned((reg321 ? wire282 : wire281)))) ?
                  reg299[(1'h0):(1'h0)] : ($unsigned(forvar316) != {reg287[(2'h2):(1'h1)]}));
            end
          else
            begin
              reg322 <= reg294;
            end
          for (forvar324 = (1'h0); (forvar324 < (3'h4)); forvar324 = (forvar324 + (1'h1)))
            begin
              reg325 = reg320;
              reg326 <= (reg288[(5'h12):(4'hc)] << (~^$unsigned((|wire280[(5'h10):(4'hd)]))));
            end
          reg327 <= (+($signed(wire281) || (((wire307 ? wire306 : reg326) ?
              wire307 : (reg313 ? reg314 : reg325)) || reg315)));
          for (forvar328 = (1'h0); (forvar328 < (2'h2)); forvar328 = (forvar328 + (1'h1)))
            begin
              reg329 <= (reg289[(1'h1):(1'h1)] >= forvar316);
              reg330 = ((wire282 ?
                  (~^$signed((-reg318))) : (+$signed($unsigned((8'hab))))) < (($signed($unsigned(reg315)) >> reg299) ?
                  wire283[(4'hc):(4'hc)] : (~({reg301} ?
                      $unsigned(reg308) : (wire307 ? reg314 : wire282)))));
              reg331 <= {$signed((-$unsigned((&reg312))))};
            end
        end
      reg332 = $unsigned((&{(8'h9c), $signed((reg312 ? reg322 : reg312))}));
      reg333 = reg315;
      reg334 = $unsigned(forvar316);
    end
  always
    @(posedge clk) begin
      if ((|wire282[(3'h5):(2'h2)]))
        begin
          if (((~|(reg294[(1'h0):(1'h0)] ?
                  (|((8'ha4) >>> (7'h43))) : (reg287 > ((7'h47) ?
                      reg290 : reg301)))) ?
              {$unsigned(($unsigned(reg289) ?
                      (reg321 ? reg329 : reg315) : reg289)),
                  ($signed((wire307 ? reg319 : reg309)) ?
                      $signed($signed(reg319)) : ((~reg305) ?
                          (reg287 << wire282) : (reg309 ?
                              reg322 : reg322)))} : (((^$signed(wire306)) <= ((&(7'h49)) - wire282)) >>> (+($signed(wire280) ?
                  (&reg301) : {reg305})))))
            begin
              reg335 <= reg290;
              reg336 = reg327[(1'h0):(1'h0)];
              reg337 <= ((((reg291[(5'h10):(2'h2)] >= $unsigned(reg288)) || ((~&reg289) ?
                          $signed((8'hb9)) : (reg299 | wire284))) ?
                      {wire282} : ($unsigned(((8'ha3) ?
                          reg305 : reg327)) && $unsigned((reg299 ?
                          (8'ha5) : reg335)))) ?
                  wire307[(3'h4):(3'h4)] : ($unsigned(((!(7'h44)) && (reg327 ?
                          reg336 : reg302))) ?
                      reg299 : $signed($signed(reg294))));
              reg338 = ($signed((^~(+$signed((8'h9e))))) < ((reg290[(2'h3):(1'h1)] + $signed(((7'h48) ?
                      reg331 : wire307))) ?
                  {((wire284 || reg302) ? {reg309, reg302} : (~|wire281)),
                      wire284[(1'h1):(1'h0)]} : $signed($unsigned((-reg309)))));
              reg339 = reg314[(3'h7):(1'h1)];
            end
          else
            begin
              reg336 = reg309[(5'h10):(1'h0)];
              reg338 = reg294[(1'h1):(1'h1)];
              reg339 = $signed((($signed((8'hbf)) ^ wire281) ?
                  $signed($signed((reg302 && reg289))) : $signed({(wire284 <= reg339),
                      $unsigned(reg294)})));
            end
        end
      else
        begin
          for (forvar335 = (1'h0); (forvar335 < (3'h4)); forvar335 = (forvar335 + (1'h1)))
            begin
              reg336 = reg288[(1'h1):(1'h0)];
              reg338 = ($unsigned($unsigned($unsigned((reg337 & wire284)))) ?
                  $signed(((-(reg338 ? (7'h4a) : reg329)) ?
                      wire284 : (reg329 ?
                          (reg339 ? reg337 : wire281) : (reg305 ?
                              (8'had) : reg335)))) : forvar335[(1'h1):(1'h0)]);
              reg339 = (-{(reg329 ? $unsigned({wire307}) : (7'h49))});
              reg340 <= (~&{($signed(((8'hbc) ? reg336 : reg305)) ?
                      $signed($signed(reg327)) : $unsigned((reg291 ?
                          wire283 : (8'ha2)))),
                  $signed($signed(wire281))});
            end
        end
    end
  assign wire341 = $signed($unsigned($signed($signed(((8'hbd) ?
                       (8'h9f) : reg322)))));
  always
    @(posedge clk) begin
      reg342 <= (wire306 ?
          (~^($signed(reg315[(2'h3):(2'h2)]) - reg326)) : $unsigned(wire306[(5'h14):(3'h5)]));
      reg343 <= (($unsigned($signed(reg340)) >= (reg321[(2'h2):(2'h2)] > reg319[(2'h3):(1'h1)])) ?
          {$signed(reg321[(2'h2):(2'h2)]),
              $signed(((reg315 ^ reg290) >> (wire307 ?
                  wire341 : reg289)))} : {$signed($signed((~(8'hb3)))),
              reg340});
      for (forvar344 = (1'h0); (forvar344 < (2'h3)); forvar344 = (forvar344 + (1'h1)))
        begin
          reg345 = reg315[(4'hf):(4'hb)];
        end
      reg346 = ($signed((((&reg337) ? $unsigned(reg294) : reg305) ?
          ($unsigned(reg345) ?
              $signed(reg287) : $signed(reg335)) : $signed(wire341[(1'h0):(1'h0)]))) <<< (|reg301[(2'h2):(1'h1)]));
      reg347 <= wire283[(4'hc):(3'h5)];
    end
  assign wire348 = $signed({reg321});
  always
    @(posedge clk) begin
      if (wire284)
        begin
          if (wire307[(3'h7):(1'h1)])
            begin
              reg349 <= (~&{$signed(($unsigned(wire306) ?
                      (8'h9d) : $unsigned(wire282)))});
              reg350 = wire284[(5'h11):(3'h6)];
            end
          else
            begin
              reg349 <= (~^(~(wire307[(2'h3):(1'h0)] ^ $signed($unsigned(reg337)))));
            end
          reg351 = reg326;
          for (forvar352 = (1'h0); (forvar352 < (1'h1)); forvar352 = (forvar352 + (1'h1)))
            begin
              reg353 = (+(7'h45));
              reg354 = reg331[(1'h1):(1'h1)];
              reg355 <= reg309;
              reg356 <= reg350;
            end
          for (forvar357 = (1'h0); (forvar357 < (3'h4)); forvar357 = (forvar357 + (1'h1)))
            begin
              reg358 = $signed($unsigned($signed($unsigned(reg337[(3'h4):(3'h4)]))));
              reg359 = $signed((reg354[(2'h3):(1'h1)] <= $signed((7'h46))));
              reg360 <= {((~&(~(reg350 + reg322))) ?
                      {reg321[(1'h0):(1'h0)]} : ((wire341 ?
                              reg359[(4'h9):(1'h0)] : reg343) ?
                          $unsigned((reg340 ~^ reg359)) : ($unsigned(wire280) ?
                              wire306[(1'h1):(1'h1)] : (wire283 ~^ reg355)))),
                  ($signed((reg353 - ((8'hbe) ? reg319 : (8'hae)))) * reg287)};
              reg361 <= ($signed(reg354) * $signed(reg315));
              reg362 <= ($signed(reg361[(2'h2):(1'h1)]) ?
                  reg301 : wire348[(4'h9):(1'h1)]);
            end
          reg363 <= {reg315};
        end
      else
        begin
          for (forvar349 = (1'h0); (forvar349 < (3'h4)); forvar349 = (forvar349 + (1'h1)))
            begin
              reg352 <= (+$signed(reg362));
              reg355 <= (({$signed($signed(reg349)), $unsigned(reg352)} ?
                  (reg299[(4'hb):(4'ha)] ?
                      reg335[(5'h13):(2'h2)] : ($unsigned(reg359) ?
                          (~reg321) : $signed(wire341))) : ((wire348[(1'h0):(1'h0)] <= reg290) ?
                      reg294 : (reg290[(2'h2):(2'h2)] ?
                          (^reg358) : (^reg353)))) >> $signed({reg331,
                  $unsigned(((8'hb8) ? reg363 : reg362))}));
              reg357 = $signed($unsigned({reg301}));
            end
          reg358 = wire280;
          reg360 <= (^~wire307);
          for (forvar361 = (1'h0); (forvar361 < (3'h4)); forvar361 = (forvar361 + (1'h1)))
            begin
              reg362 <= {($unsigned(($unsigned(reg299) <= reg351[(3'h4):(1'h1)])) ?
                      wire306[(4'he):(4'h9)] : ((reg353[(3'h4):(2'h2)] + $signed(wire348)) ~^ reg337[(4'h8):(3'h6)]))};
              reg363 <= $signed(reg351);
              reg364 <= ((((|(reg319 + reg287)) ?
                      ({reg358} ?
                          reg355[(4'hb):(3'h5)] : (~^wire348)) : reg361[(3'h6):(1'h1)]) ?
                  {{$signed(reg289)},
                      (-reg356[(4'he):(4'hc)])} : reg315) < $signed(reg319[(2'h2):(2'h2)]));
              reg365 = ({reg356,
                      (reg358[(4'hb):(3'h6)] ?
                          $unsigned(reg302[(2'h2):(2'h2)]) : ((-reg294) ?
                              $signed(reg331) : $unsigned(reg343)))} ?
                  ($unsigned({$unsigned(reg327)}) + ($unsigned((wire284 * reg309)) >>> $unsigned({reg362}))) : ((^$signed((&reg364))) ?
                      $unsigned(((!(8'hac)) & {wire348,
                          forvar349})) : (8'ha0)));
            end
        end
      if ((reg314 ? reg349[(4'h8):(1'h0)] : reg357))
        begin
          reg366 = ((wire306 <= (reg342[(1'h1):(1'h0)] > reg299[(2'h3):(1'h0)])) ^~ ((reg358[(2'h3):(2'h2)] ~^ reg305[(4'h9):(1'h0)]) || ((+{reg302}) | $signed((8'ha4)))));
          reg367 = reg302[(4'h9):(3'h4)];
        end
      else
        begin
          if (wire307[(4'h9):(2'h2)])
            begin
              reg368 <= (({$unsigned((-forvar349)),
                  (reg327 ?
                      $unsigned(reg301) : ((7'h47) ?
                          reg340 : reg357))} || (-reg302[(4'h9):(3'h6)])) || (~&{($unsigned(reg349) ?
                      (reg349 || reg342) : ((8'ha0) ? reg327 : reg357)),
                  (+wire284[(4'h8):(2'h2)])}));
              reg369 <= $signed((^forvar349[(4'h9):(4'h8)]));
            end
          else
            begin
              reg368 <= $unsigned(($unsigned(((~&wire281) || forvar352)) * (((reg294 ~^ (8'h9e)) ?
                  (~(8'ha5)) : reg352[(3'h7):(2'h3)]) + (reg342[(3'h5):(1'h0)] >>> (+reg294)))));
              reg369 <= reg357;
              reg370 <= (wire306[(3'h7):(3'h6)] ? (reg349 ^ (7'h44)) : reg368);
              reg371 = reg315[(2'h2):(2'h2)];
              reg372 = (&reg343);
            end
          reg373 <= (reg343 ?
              wire307[(4'hb):(3'h5)] : (&$unsigned({(reg287 ? (8'hbe) : reg321),
                  $unsigned(reg366)})));
        end
      reg374 = ($unsigned(((~|wire282) ~^ reg329[(3'h6):(2'h2)])) != (wire284 ?
          $unsigned(reg335) : (forvar349 ?
              $unsigned($signed(reg370)) : ($signed(reg370) > (reg362 ?
                  reg326 : reg372)))));
    end
  always
    @(posedge clk) begin
      if ($unsigned((|$unsigned((~|(!reg362))))))
        begin
          reg375 = ((^~(($unsigned(wire341) ? ((8'hae) != reg290) : (!reg305)) ?
              $unsigned({reg349}) : wire307[(2'h2):(2'h2)])) ^ reg287[(3'h5):(3'h4)]);
          for (forvar376 = (1'h0); (forvar376 < (2'h2)); forvar376 = (forvar376 + (1'h1)))
            begin
              reg377 = {reg315[(2'h2):(1'h1)]};
              reg378 <= (reg321[(2'h2):(2'h2)] >>> $signed($unsigned(reg301[(2'h2):(2'h2)])));
              reg379 = $signed(reg363[(4'hb):(4'ha)]);
              reg380 = reg289;
              reg381 <= $signed(((8'hbb) <= ($signed($unsigned(wire307)) ?
                  reg321[(3'h4):(3'h4)] : $unsigned((reg377 & (8'ha4))))));
            end
        end
      else
        begin
          reg376 <= reg352;
          reg377 = $signed((+{reg302}));
          reg379 = ($unsigned($unsigned($unsigned((wire306 ^ reg381)))) ?
              reg290 : (reg314[(3'h7):(3'h4)] ?
                  (^(~^(!wire341))) : {($unsigned(reg375) <<< $signed(reg342))}));
        end
      for (forvar382 = (1'h0); (forvar382 < (2'h2)); forvar382 = (forvar382 + (1'h1)))
        begin
          reg383 = (!(8'ha2));
        end
      for (forvar384 = (1'h0); (forvar384 < (3'h4)); forvar384 = (forvar384 + (1'h1)))
        begin
          if ($signed(((!$signed(forvar376[(4'h8):(1'h1)])) ?
              $signed(reg315[(4'ha):(4'h8)]) : ($unsigned((reg337 * reg340)) | (^$signed(wire281))))))
            begin
              reg385 <= (^~(-$signed(reg331)));
              reg386 <= $signed($unsigned($unsigned(($unsigned((8'haa)) ?
                  (+(7'h41)) : $signed((8'ha2))))));
              reg387 <= reg347[(1'h1):(1'h0)];
              reg388 <= {$signed($unsigned($unsigned((wire348 <= reg386)))),
                  {reg373, ($signed($unsigned((7'h41))) && reg301)}};
            end
          else
            begin
              reg389 = (~^(8'ha3));
              reg390 = ($unsigned(reg362[(3'h4):(3'h4)]) ?
                  $signed($unsigned(({reg340} == (^wire281)))) : $signed(($signed((reg361 ^~ reg378)) ?
                      reg360 : reg287)));
              reg391 = {((({reg321, reg383} || $unsigned(wire282)) ?
                      $unsigned(reg373) : wire307[(4'hb):(4'h9)]) ~^ reg389)};
            end
        end
    end
  assign wire392 = (reg329[(2'h2):(2'h2)] ?
                       (reg376 ^ ((^~(-reg294)) == (reg349[(1'h1):(1'h0)] < (reg290 ?
                           wire280 : reg305)))) : reg288[(5'h13):(5'h13)]);
  assign wire393 = (({$signed(reg289[(3'h5):(1'h1)]), $unsigned({(8'hb9)})} ?
                       (({reg302, reg343} >> (^(8'hbb))) ?
                           ($unsigned(wire306) ?
                               $unsigned(reg356) : (&reg373)) : {(^~reg373)}) : reg361[(3'h6):(1'h1)]) ^ {($signed({wire280}) ?
                           ($unsigned((8'hbe)) && (reg301 ?
                               (8'hb0) : (8'had))) : (reg343 ?
                               reg387[(4'hd):(2'h3)] : $unsigned(reg347)))});
  module394 #() modinst427 (wire426, clk, reg290, reg319, reg322, wire392);
  module428 #() modinst623 (.wire430(wire282), .clk(clk), .wire431(reg387), .wire432(reg368), .wire433(reg299), .wire429(wire426), .y(wire622));
  assign wire624 = (wire306 <<< (^{reg347[(1'h0):(1'h0)],
                       $unsigned($unsigned((8'ha3)))}));
  always
    @(posedge clk) begin
      reg625 = (-$unsigned({(wire392[(4'he):(4'ha)] > (reg329 ?
              reg386 : reg385))}));
      reg626 = (($signed($unsigned($signed(wire393))) ?
          wire348 : $signed((8'ha0))) >= (($unsigned((8'haf)) ^~ $unsigned({wire392})) >> $unsigned((reg305[(2'h2):(2'h2)] ?
          reg327 : (+reg309)))));
      for (forvar627 = (1'h0); (forvar627 < (1'h0)); forvar627 = (forvar627 + (1'h1)))
        begin
          reg628 = $signed({(+$signed(wire284))});
          reg629 <= (wire283[(4'h8):(3'h5)] ?
              (reg305 & (reg289[(3'h6):(2'h3)] >= (~&(8'ha4)))) : ($unsigned((~|(reg337 ?
                      wire284 : wire341))) ?
                  ((~^reg376) ?
                      ((8'hb3) ?
                          reg363[(3'h7):(3'h7)] : $signed(reg347)) : wire307) : reg342[(1'h0):(1'h0)]));
        end
    end
  assign wire630 = $unsigned($unsigned($unsigned((~reg301[(4'h8):(3'h6)]))));
  always
    @(posedge clk) begin
      if (($signed(reg291[(1'h1):(1'h1)]) >>> ($signed($unsigned($unsigned(reg309))) ?
          $signed(((-(8'hb9)) ?
              $unsigned(reg305) : (reg361 < reg356))) : wire392[(4'ha):(4'h8)])))
        begin
          reg631 <= reg331;
          reg632 <= reg322[(5'h13):(4'ha)];
        end
      else
        begin
          reg631 <= reg355[(4'ha):(3'h5)];
          reg632 <= $signed({reg370[(1'h1):(1'h1)], $unsigned(reg378)});
        end
      for (forvar633 = (1'h0); (forvar633 < (1'h0)); forvar633 = (forvar633 + (1'h1)))
        begin
          reg634 <= $unsigned((+($signed((wire426 != wire284)) ?
              reg387[(4'h8):(3'h7)] : ($signed(reg331) ?
                  (reg349 << reg326) : reg363[(3'h4):(2'h2)]))));
          for (forvar635 = (1'h0); (forvar635 < (2'h2)); forvar635 = (forvar635 + (1'h1)))
            begin
              reg636 = {reg337,
                  (~|(reg373 >= $signed((reg331 ? (8'hb2) : reg329))))};
              reg637 <= reg287[(3'h5):(1'h1)];
              reg638 <= {$unsigned({($signed(wire283) ~^ (!wire307))})};
            end
          reg639 = (reg314[(2'h3):(2'h2)] ?
              $signed(wire284[(3'h4):(1'h0)]) : (^~$signed((reg343[(3'h5):(1'h0)] | (reg631 <<< (8'hba))))));
          for (forvar640 = (1'h0); (forvar640 < (2'h3)); forvar640 = (forvar640 + (1'h1)))
            begin
              reg641 <= reg342;
              reg642 <= reg302[(4'hd):(3'h5)];
            end
          for (forvar643 = (1'h0); (forvar643 < (1'h1)); forvar643 = (forvar643 + (1'h1)))
            begin
              reg644 = $unsigned((~&(|wire622[(2'h2):(1'h1)])));
              reg645 <= (^~reg636);
              reg646 <= reg381[(4'hf):(4'hc)];
              reg647 = (reg309 || reg364);
              reg648 = reg376;
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module428
#(parameter param621 = ({((~^((7'h43) + (8'haf))) | ((8'haa) ? ((8'hbf) >= (8'ha4)) : (~|(7'h47)))), ((^(~&(8'ha1))) || ((|(8'ha9)) ? (8'hbe) : (&(7'h40))))} ? (((((8'hb1) ? (8'hb9) : (8'haf)) ? (8'hb0) : (8'hb9)) ? (((8'ha9) == (8'hb4)) >>> (^~(8'ha3))) : {((8'hb1) ? (7'h48) : (8'ha8)), {(7'h41)}}) ? ((+(~^(7'h49))) >> (((8'h9d) > (7'h40)) ? ((7'h42) ? (8'hb1) : (8'hb1)) : ((8'hab) ? (8'had) : (8'hb5)))) : (({(8'ha4), (8'haa)} > {(8'hbe), (7'h4a)}) ? (^{(8'hb4)}) : (&{(8'hac)}))) : (8'ha4)))
(y, clk, wire433, wire432, wire431, wire430, wire429);
  output wire [(32'h9db):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire433;
  input wire [(3'h7):(1'h0)] wire432;
  input wire [(5'h10):(1'h0)] wire431;
  input wire [(4'hb):(1'h0)] wire430;
  input wire [(3'h4):(1'h0)] wire429;
  wire signed [(2'h3):(1'h0)] wire567;
  wire signed [(4'h9):(1'h0)] wire566;
  wire signed [(5'h14):(1'h0)] wire465;
  wire signed [(4'h8):(1'h0)] wire464;
  wire [(4'h8):(1'h0)] wire435;
  wire signed [(5'h11):(1'h0)] wire434;
  reg [(4'h8):(1'h0)] reg620 = (1'h0);
  reg [(5'h14):(1'h0)] reg619 = (1'h0);
  reg [(3'h5):(1'h0)] reg613 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg612 = (1'h0);
  reg [(5'h18):(1'h0)] reg611 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg610 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg608 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg607 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg604 = (1'h0);
  reg [(5'h15):(1'h0)] reg603 = (1'h0);
  reg [(5'h18):(1'h0)] reg600 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg599 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg594 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg592 = (1'h0);
  reg [(5'h15):(1'h0)] reg589 = (1'h0);
  reg [(5'h14):(1'h0)] reg588 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg586 = (1'h0);
  reg [(4'h8):(1'h0)] reg584 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg582 = (1'h0);
  reg [(4'hf):(1'h0)] reg578 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg575 = (1'h0);
  reg [(3'h6):(1'h0)] reg571 = (1'h0);
  reg [(5'h12):(1'h0)] reg563 = (1'h0);
  reg signed [(4'he):(1'h0)] reg560 = (1'h0);
  reg [(4'h8):(1'h0)] reg557 = (1'h0);
  reg [(3'h6):(1'h0)] reg555 = (1'h0);
  reg [(5'h15):(1'h0)] reg553 = (1'h0);
  reg [(4'he):(1'h0)] reg552 = (1'h0);
  reg [(4'ha):(1'h0)] reg549 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg547 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg544 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg542 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg540 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg519 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg533 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg532 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg531 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg529 = (1'h0);
  reg [(4'hb):(1'h0)] reg528 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg527 = (1'h0);
  reg [(5'h10):(1'h0)] reg526 = (1'h0);
  reg [(4'hb):(1'h0)] reg525 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg520 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg518 = (1'h0);
  reg [(5'h17):(1'h0)] reg512 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg503 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg508 = (1'h0);
  reg [(3'h7):(1'h0)] reg506 = (1'h0);
  reg [(5'h14):(1'h0)] reg501 = (1'h0);
  reg [(5'h10):(1'h0)] reg498 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg497 = (1'h0);
  reg [(4'hf):(1'h0)] reg496 = (1'h0);
  reg [(4'hf):(1'h0)] reg495 = (1'h0);
  reg [(5'h18):(1'h0)] reg494 = (1'h0);
  reg [(4'he):(1'h0)] reg493 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg491 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg490 = (1'h0);
  reg [(5'h15):(1'h0)] reg488 = (1'h0);
  reg [(5'h12):(1'h0)] reg486 = (1'h0);
  reg [(5'h11):(1'h0)] reg485 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg481 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg477 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg474 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg472 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg471 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg469 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg461 = (1'h0);
  reg [(5'h16):(1'h0)] reg459 = (1'h0);
  reg [(5'h18):(1'h0)] reg458 = (1'h0);
  reg signed [(4'he):(1'h0)] reg457 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg451 = (1'h0);
  reg [(2'h3):(1'h0)] reg450 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg446 = (1'h0);
  reg [(4'he):(1'h0)] reg442 = (1'h0);
  reg [(4'h8):(1'h0)] reg440 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg439 = (1'h0);
  reg [(4'hd):(1'h0)] reg438 = (1'h0);
  reg [(3'h5):(1'h0)] reg437 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg618 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg617 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg616 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg615 = (1'h0);
  reg [(5'h10):(1'h0)] reg614 = (1'h0);
  reg signed [(4'he):(1'h0)] reg609 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg606 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg605 = (1'h0);
  reg [(3'h4):(1'h0)] reg602 = (1'h0);
  reg [(4'h8):(1'h0)] reg601 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg598 = (1'h0);
  reg [(4'h9):(1'h0)] reg597 = (1'h0);
  reg [(3'h5):(1'h0)] reg596 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg593 = (1'h0);
  reg signed [(4'he):(1'h0)] reg591 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg590 = (1'h0);
  reg [(4'ha):(1'h0)] reg587 = (1'h0);
  reg [(4'h8):(1'h0)] reg585 = (1'h0);
  reg [(4'he):(1'h0)] reg583 = (1'h0);
  reg [(3'h6):(1'h0)] reg581 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar580 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg579 = (1'h0);
  reg [(5'h13):(1'h0)] reg577 = (1'h0);
  reg [(5'h13):(1'h0)] reg576 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg574 = (1'h0);
  reg [(5'h16):(1'h0)] reg573 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg572 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg570 = (1'h0);
  reg [(4'h9):(1'h0)] forvar569 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar568 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg565 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg564 = (1'h0);
  reg [(2'h3):(1'h0)] forvar562 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg561 = (1'h0);
  reg [(3'h7):(1'h0)] reg559 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg558 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg556 = (1'h0);
  reg [(5'h14):(1'h0)] reg554 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar551 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar550 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg548 = (1'h0);
  reg [(4'ha):(1'h0)] reg546 = (1'h0);
  reg [(4'hd):(1'h0)] forvar545 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg543 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg541 = (1'h0);
  reg [(4'ha):(1'h0)] reg539 = (1'h0);
  reg [(4'ha):(1'h0)] reg538 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg537 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar536 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar526 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar518 = (1'h0);
  reg [(4'hd):(1'h0)] reg535 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg534 = (1'h0);
  reg [(4'hf):(1'h0)] reg530 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg524 = (1'h0);
  reg [(3'h6):(1'h0)] reg523 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg522 = (1'h0);
  reg [(5'h15):(1'h0)] reg521 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar519 = (1'h0);
  reg [(3'h6):(1'h0)] reg517 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg516 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg515 = (1'h0);
  reg [(4'hf):(1'h0)] reg514 = (1'h0);
  reg [(4'h8):(1'h0)] reg513 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar511 = (1'h0);
  reg signed [(4'he):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar505 = (1'h0);
  reg [(3'h5):(1'h0)] reg507 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg505 = (1'h0);
  reg [(5'h13):(1'h0)] reg504 = (1'h0);
  reg [(2'h3):(1'h0)] forvar503 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg502 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg500 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg499 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg492 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar481 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar479 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg489 = (1'h0);
  reg [(5'h10):(1'h0)] reg487 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg484 = (1'h0);
  reg [(5'h16):(1'h0)] reg483 = (1'h0);
  reg [(3'h5):(1'h0)] reg482 = (1'h0);
  reg [(5'h13):(1'h0)] reg480 = (1'h0);
  reg [(2'h3):(1'h0)] reg479 = (1'h0);
  reg [(5'h18):(1'h0)] forvar478 = (1'h0);
  reg [(5'h16):(1'h0)] reg476 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg475 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar470 = (1'h0);
  reg [(5'h16):(1'h0)] reg473 = (1'h0);
  reg [(4'he):(1'h0)] reg470 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg468 = (1'h0);
  reg [(3'h7):(1'h0)] reg467 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg466 = (1'h0);
  reg [(4'h8):(1'h0)] reg463 = (1'h0);
  reg [(5'h14):(1'h0)] reg462 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg460 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg456 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg455 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg454 = (1'h0);
  reg [(5'h17):(1'h0)] reg453 = (1'h0);
  reg [(3'h4):(1'h0)] reg452 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg449 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg448 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar447 = (1'h0);
  reg [(3'h6):(1'h0)] reg445 = (1'h0);
  reg [(3'h5):(1'h0)] reg444 = (1'h0);
  reg [(4'hb):(1'h0)] reg443 = (1'h0);
  reg [(4'he):(1'h0)] forvar437 = (1'h0);
  reg [(3'h5):(1'h0)] reg441 = (1'h0);
  reg [(2'h2):(1'h0)] reg436 = (1'h0);
  assign y = {wire567,
                 wire566,
                 wire465,
                 wire464,
                 wire435,
                 wire434,
                 reg620,
                 reg619,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 reg608,
                 reg607,
                 reg604,
                 reg603,
                 reg600,
                 reg599,
                 reg594,
                 reg592,
                 reg589,
                 reg588,
                 reg586,
                 reg584,
                 reg582,
                 reg578,
                 reg575,
                 reg571,
                 reg563,
                 reg560,
                 reg557,
                 reg555,
                 reg553,
                 reg552,
                 reg549,
                 reg547,
                 reg544,
                 reg542,
                 reg540,
                 reg519,
                 reg533,
                 reg532,
                 reg531,
                 reg529,
                 reg528,
                 reg527,
                 reg526,
                 reg525,
                 reg520,
                 reg518,
                 reg512,
                 reg510,
                 reg503,
                 reg508,
                 reg506,
                 reg501,
                 reg498,
                 reg497,
                 reg496,
                 reg495,
                 reg494,
                 reg493,
                 reg491,
                 reg490,
                 reg488,
                 reg486,
                 reg485,
                 reg481,
                 reg477,
                 reg474,
                 reg472,
                 reg471,
                 reg469,
                 reg461,
                 reg459,
                 reg458,
                 reg457,
                 reg451,
                 reg450,
                 reg446,
                 reg442,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg618,
                 reg617,
                 reg616,
                 reg615,
                 reg614,
                 reg609,
                 reg606,
                 reg605,
                 reg602,
                 reg601,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 reg593,
                 reg591,
                 reg590,
                 reg587,
                 reg585,
                 reg583,
                 reg581,
                 forvar580,
                 reg579,
                 reg577,
                 reg576,
                 reg574,
                 reg573,
                 reg572,
                 reg570,
                 forvar569,
                 forvar568,
                 reg565,
                 reg564,
                 forvar562,
                 reg561,
                 reg559,
                 reg558,
                 reg556,
                 reg554,
                 forvar551,
                 forvar550,
                 reg548,
                 reg546,
                 forvar545,
                 reg543,
                 reg541,
                 reg539,
                 reg538,
                 reg537,
                 forvar536,
                 forvar526,
                 forvar518,
                 reg535,
                 reg534,
                 reg530,
                 reg524,
                 reg523,
                 reg522,
                 reg521,
                 forvar519,
                 reg517,
                 reg516,
                 reg515,
                 reg514,
                 reg513,
                 forvar511,
                 reg509,
                 forvar505,
                 reg507,
                 reg505,
                 reg504,
                 forvar503,
                 reg502,
                 reg500,
                 reg499,
                 reg492,
                 forvar481,
                 forvar479,
                 reg478,
                 reg489,
                 reg487,
                 reg484,
                 reg483,
                 reg482,
                 reg480,
                 reg479,
                 forvar478,
                 reg476,
                 reg475,
                 forvar470,
                 reg473,
                 reg470,
                 reg468,
                 reg467,
                 reg466,
                 reg463,
                 reg462,
                 reg460,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg449,
                 reg448,
                 forvar447,
                 reg445,
                 reg444,
                 reg443,
                 forvar437,
                 reg441,
                 reg436,
                 (1'h0)};
  assign wire434 = $unsigned(({(wire429 ?
                           (wire429 ? wire431 : wire433) : $signed(wire430)),
                       $signed(wire433)} * $unsigned(wire433[(2'h3):(2'h3)])));
  assign wire435 = wire432;
  always
    @(posedge clk) begin
      reg436 = wire432[(2'h3):(2'h2)];
      if ({(8'haf)})
        begin
          if ($unsigned(($signed(((wire435 ? wire432 : reg436) + (wire433 ?
                  wire430 : wire430))) ?
              (^~$unsigned(wire430[(3'h6):(3'h5)])) : $signed(wire431))))
            begin
              reg437 <= ($signed(wire430) ^~ {wire434[(2'h2):(1'h0)],
                  $signed(wire429)});
              reg438 <= {wire433[(4'ha):(2'h3)], $signed($signed(wire432))};
              reg439 <= (wire433[(1'h0):(1'h0)] * wire433);
              reg440 <= wire435;
            end
          else
            begin
              reg437 <= wire433;
              reg438 <= {$unsigned(reg436[(1'h1):(1'h1)])};
              reg439 <= $unsigned(({wire430, reg439[(4'hc):(3'h7)]} ?
                  (~(~(wire433 - reg437))) : (wire430 ?
                      ((~^reg438) ?
                          $unsigned(wire435) : $unsigned(wire431)) : (-$unsigned(wire431)))));
            end
          reg441 = $signed($signed($unsigned(wire432)));
        end
      else
        begin
          for (forvar437 = (1'h0); (forvar437 < (2'h2)); forvar437 = (forvar437 + (1'h1)))
            begin
              reg438 <= ((~^(($signed(wire430) ?
                          (reg440 >> forvar437) : (wire429 < wire433)) ?
                      wire433[(4'hd):(1'h1)] : reg437)) ?
                  ({(^~reg440)} & $unsigned((|reg436))) : ($signed($signed({reg437})) > ($unsigned((~wire434)) & $signed(wire432[(3'h4):(1'h1)]))));
              reg439 <= reg441[(2'h2):(1'h1)];
            end
          if (reg441[(1'h1):(1'h0)])
            begin
              reg441 = $signed((&wire430));
            end
          else
            begin
              reg441 = reg436;
              reg442 <= reg438[(3'h5):(2'h2)];
              reg443 = $unsigned($unsigned(((+reg436) >>> $unsigned((wire435 ?
                  wire431 : reg436)))));
              reg444 = ((-reg439) ?
                  wire429[(3'h4):(1'h1)] : (reg443[(3'h4):(1'h0)] ?
                      reg441 : $signed((&$unsigned(wire432)))));
            end
          if (($unsigned($unsigned(reg437[(3'h4):(2'h2)])) ?
              $unsigned(reg438[(1'h1):(1'h0)]) : ($unsigned((reg437[(3'h4):(1'h1)] - (^wire433))) & (((reg443 ?
                          wire433 : wire431) ?
                      $unsigned(reg438) : (~&reg444)) ?
                  ($unsigned(reg444) <<< $unsigned(reg439)) : {(~wire434)}))))
            begin
              reg445 = $signed({((^~reg443) || ((reg439 != wire433) ?
                      wire434 : $signed(wire435))),
                  wire430});
            end
          else
            begin
              reg446 <= (^~(8'hbe));
            end
          for (forvar447 = (1'h0); (forvar447 < (1'h1)); forvar447 = (forvar447 + (1'h1)))
            begin
              reg448 = $signed($signed((-{wire429, reg436[(1'h1):(1'h1)]})));
              reg449 = $signed({((wire429 ?
                      ((7'h43) & (8'h9d)) : $signed(reg436)) << reg437),
                  $unsigned((|(reg443 << reg436)))});
              reg450 <= wire430;
              reg451 <= reg443;
            end
        end
      reg452 = $unsigned(($signed(wire435) ?
          ((wire435 ? (&reg451) : (reg449 >> reg449)) ?
              (reg436 >>> $unsigned(wire431)) : reg445) : {{(reg441 | reg444)}}));
      reg453 = $signed((~|(reg436[(1'h1):(1'h1)] ?
          ((wire430 + reg451) || (reg449 ?
              forvar437 : forvar447)) : (((8'haf) >= reg439) ?
              $signed(reg448) : (8'ha7)))));
    end
  always
    @(posedge clk) begin
      if ($unsigned((8'ha2)))
        begin
          reg454 = wire433[(3'h7):(3'h6)];
          reg455 = $signed(reg438);
          if ($signed($unsigned(reg451[(3'h4):(2'h3)])))
            begin
              reg456 = wire434;
            end
          else
            begin
              reg457 <= $signed($signed((reg451 ~^ {reg442})));
              reg458 <= reg450[(1'h1):(1'h1)];
              reg459 <= $signed((((|$unsigned(reg457)) * ($unsigned((8'hbc)) & $signed((8'h9f)))) ?
                  $signed(wire429) : ((wire431 ?
                          (reg438 == (8'ha9)) : $unsigned(reg438)) ?
                      $signed(reg446) : $unsigned({wire431, reg454}))));
            end
          reg460 = (~&({(((7'h47) ?
                  wire430 : wire434) ~^ reg456[(4'h9):(3'h7)]),
              reg457[(4'h8):(1'h1)]} ^ ($unsigned((^~(7'h40))) || $unsigned($signed(reg456)))));
        end
      else
        begin
          if ($signed(wire432[(3'h6):(3'h6)]))
            begin
              reg454 = ((7'h47) ? reg454 : (^~{reg446}));
            end
          else
            begin
              reg454 = ($signed(reg439[(2'h2):(1'h1)]) ?
                  $signed(($signed((reg456 <= reg440)) < (&(reg451 ^~ wire433)))) : $unsigned($signed((^~(wire430 ?
                      wire432 : (7'h42))))));
              reg455 = {(((~&$signed(reg460)) << ({wire430,
                          reg451} ^~ (reg458 << wire434))) ?
                      reg439[(1'h1):(1'h0)] : ((+wire431) ?
                          $signed($unsigned(reg456)) : {$signed(reg456)}))};
            end
          if ({reg446})
            begin
              reg456 = $unsigned($unsigned({$signed(reg458[(5'h15):(3'h5)])}));
              reg457 <= (reg438 ?
                  (+((&$signed(reg450)) ?
                      ($signed(reg440) >> (7'h4a)) : (^(wire432 ?
                          reg456 : reg455)))) : {reg442[(4'hb):(3'h6)],
                      (~&wire433[(3'h4):(2'h2)])});
              reg460 = (wire430[(3'h4):(1'h1)] + {($unsigned($signed(wire430)) ?
                      reg459 : reg455[(4'hb):(2'h2)]),
                  $unsigned($unsigned(reg446))});
              reg461 <= (((!$signed(reg454)) ?
                  wire434 : {reg439,
                      $signed($signed(reg439))}) > $signed(reg458[(4'ha):(2'h3)]));
            end
          else
            begin
              reg456 = $unsigned($unsigned({{{reg438}, (reg459 >> (8'hb6))}}));
              reg457 <= $signed(($unsigned(({reg458,
                  reg437} ^~ (8'had))) & reg459));
              reg460 = ((~reg460[(2'h3):(2'h2)]) | (&(reg450[(2'h2):(1'h1)] + $unsigned(reg454))));
              reg462 = $unsigned((8'hb1));
            end
          reg463 = reg462[(3'h6):(1'h0)];
        end
    end
  assign wire464 = {$unsigned($signed($signed(((7'h41) + (8'ha6))))),
                       (wire430 ~^ ({(|reg458), (reg442 > reg458)} ?
                           reg457 : {reg451[(2'h3):(1'h1)]}))};
  assign wire465 = (^(wire434 ?
                       $unsigned(wire435[(2'h2):(1'h1)]) : {wire430[(4'h9):(1'h1)]}));
  always
    @(posedge clk) begin
      if (((~&{(!{wire431}), reg437}) ?
          wire429[(1'h1):(1'h1)] : ($unsigned((~|reg438)) * (((reg450 + wire433) << reg438[(4'hd):(3'h4)]) ?
              reg461[(4'hc):(1'h1)] : $signed((&(8'hb9)))))))
        begin
          if ($unsigned((8'ha6)))
            begin
              reg466 = (~({wire431[(4'ha):(3'h7)]} ?
                  (reg450 ^ ($signed(wire435) * wire434[(5'h10):(2'h3)])) : $signed({(^~wire433)})));
              reg467 = $signed(wire431);
              reg468 = {reg466};
            end
          else
            begin
              reg466 = ((^~((|reg461) ~^ ((reg467 ^~ reg466) ?
                      (wire464 ? (7'h44) : wire430) : (wire429 * reg446)))) ?
                  $unsigned((wire429[(3'h4):(1'h0)] ?
                      reg446[(3'h5):(3'h4)] : (wire431 ?
                          (^~reg466) : wire431))) : ((reg466 ?
                          $unsigned({reg468, reg442}) : reg446[(3'h7):(2'h3)]) ?
                      wire432 : (8'ha6)));
              reg467 = $signed((-reg437));
              reg469 <= ((((!reg440[(1'h0):(1'h0)]) ?
                          reg438 : ((!wire464) * $unsigned(reg467))) ?
                      {(wire429 >> $unsigned((8'ha4)))} : reg437) ?
                  (8'hbd) : {$unsigned($signed(((8'ha6) ? reg440 : reg442))),
                      (reg437 ?
                          $unsigned((wire432 >>> (8'hb0))) : (^(wire433 && wire429)))});
            end
          reg470 = (wire434[(3'h6):(1'h1)] ?
              {({(wire430 + wire431),
                      (wire432 || (8'ha0))} * (^reg459[(4'hd):(1'h1)]))} : reg451[(2'h2):(1'h0)]);
          reg471 <= reg461;
          reg472 <= ((|wire435[(2'h3):(2'h3)]) >> reg457);
          reg473 = $unsigned((-reg461));
        end
      else
        begin
          reg469 <= wire434[(3'h6):(3'h4)];
          for (forvar470 = (1'h0); (forvar470 < (1'h0)); forvar470 = (forvar470 + (1'h1)))
            begin
              reg473 = ($unsigned((reg439 ?
                      ({(8'hb0), reg472} ^~ ((8'hb9) != reg472)) : reg467)) ?
                  ($unsigned($signed((^~(8'h9d)))) ?
                      (-$unsigned($signed(wire433))) : $unsigned({(8'ha2)})) : ((7'h43) << ((~|reg438) ^ {reg467,
                      (reg440 && reg437)})));
              reg474 <= ($signed((~|(~(-wire464)))) ?
                  (reg459[(5'h12):(4'h8)] == {wire434[(4'hd):(4'h9)],
                      (~|reg440[(3'h5):(2'h3)])}) : ($signed((~$unsigned(wire435))) ?
                      (7'h46) : ($unsigned((reg450 > reg458)) ?
                          reg461 : $signed(reg440[(3'h5):(1'h0)]))));
            end
          if ((8'hb4))
            begin
              reg475 = reg470[(3'h4):(2'h2)];
            end
          else
            begin
              reg475 = reg473;
              reg476 = {$signed(wire433)};
            end
          reg477 <= (-reg469);
        end
      if (reg461[(4'hd):(3'h4)])
        begin
          for (forvar478 = (1'h0); (forvar478 < (2'h3)); forvar478 = (forvar478 + (1'h1)))
            begin
              reg479 = wire465;
              reg480 = $signed($unsigned($unsigned((^reg473[(5'h10):(4'hb)]))));
              reg481 <= $signed((wire429 ? {wire464} : reg480[(5'h12):(4'hf)]));
              reg482 = $unsigned(reg474[(5'h11):(4'hb)]);
              reg483 = (~^$unsigned((+wire429)));
            end
          reg484 = reg479[(2'h2):(2'h2)];
          if (((reg437 ?
                  {reg484, (8'ha8)} : (wire465[(4'ha):(1'h1)] ?
                      reg477[(4'h9):(4'h8)] : (((8'hb2) << reg442) <= (reg474 >> reg439)))) ?
              $unsigned((((!reg450) ?
                  $signed(wire465) : {reg482}) ~^ $signed(reg481[(4'h8):(3'h6)]))) : reg482))
            begin
              reg485 <= (wire429[(1'h0):(1'h0)] ?
                  $unsigned((~^wire429)) : reg457);
              reg486 <= ({reg458,
                  (($unsigned((8'ha7)) != (reg482 || reg473)) ?
                      $signed((reg480 ?
                          reg468 : (8'hb8))) : reg442[(3'h5):(3'h5)])} >>> $signed(reg481[(4'hb):(3'h5)]));
            end
          else
            begin
              reg487 = (+reg483);
              reg488 <= ($unsigned(wire434) ?
                  (reg440[(4'h8):(3'h6)] ?
                      (~^($signed(reg471) < (reg476 ?
                          reg438 : (8'hb4)))) : (((wire433 ?
                                  (7'h47) : wire432) ?
                              (reg457 * (8'ha8)) : (~^reg457)) ?
                          reg451[(3'h5):(3'h5)] : (8'hae))) : $signed((wire429[(1'h1):(1'h0)] ?
                      wire435[(3'h5):(1'h0)] : ($unsigned(wire429) ^ {wire464,
                          reg483}))));
              reg489 = {reg483[(5'h15):(5'h14)]};
            end
          reg490 <= reg440;
        end
      else
        begin
          reg478 = (&((^($signed(reg457) ? forvar478[(4'hd):(3'h4)] : reg450)) ?
              wire465[(5'h13):(5'h12)] : $unsigned(((wire465 ?
                  wire430 : (7'h43)) >>> reg490))));
          for (forvar479 = (1'h0); (forvar479 < (2'h3)); forvar479 = (forvar479 + (1'h1)))
            begin
              reg480 = reg438[(4'hb):(3'h4)];
            end
          for (forvar481 = (1'h0); (forvar481 < (2'h3)); forvar481 = (forvar481 + (1'h1)))
            begin
              reg485 <= (&(($unsigned($unsigned(reg481)) ?
                  $unsigned((reg468 ?
                      wire435 : reg476)) : $unsigned((+reg476))) || (~$signed($unsigned(reg470)))));
              reg487 = ((~^$unsigned(((reg450 >> reg490) & (7'h44)))) ?
                  {(reg483 ?
                          ($unsigned(reg442) ~^ {wire429}) : (!$signed(reg472))),
                      $unsigned({(reg459 ~^ wire432),
                          (^reg477)})} : $unsigned(reg473[(5'h11):(4'he)]));
              reg488 <= $unsigned($unsigned(reg438));
            end
          if ($unsigned($unsigned(($unsigned({reg438}) ?
              ((reg470 << (8'hbf)) == (!reg470)) : (reg457 == $unsigned(forvar470))))))
            begin
              reg490 <= (reg478[(3'h5):(3'h4)] ?
                  reg437[(2'h2):(2'h2)] : ($unsigned({(~&wire433),
                      (^reg486)}) < wire431[(3'h5):(1'h1)]));
              reg491 <= $unsigned($unsigned($unsigned($unsigned($unsigned(reg472)))));
              reg492 = (^(~&reg439));
              reg493 <= (~|reg451);
              reg494 <= {($unsigned((((8'hbb) > reg478) <<< (reg485 ?
                      reg438 : wire435))) ^ $signed(reg459))};
            end
          else
            begin
              reg489 = forvar470[(4'hb):(2'h2)];
              reg492 = $unsigned(reg451[(3'h4):(3'h4)]);
              reg493 <= forvar478[(3'h5):(1'h0)];
              reg494 <= {(^reg481[(3'h4):(2'h2)])};
            end
        end
    end
  always
    @(posedge clk) begin
      if ($signed({(wire430[(2'h3):(2'h2)] ?
              wire465[(4'hb):(4'h8)] : $signed({(8'hbb), reg494})),
          reg457}))
        begin
          reg495 <= reg446;
          reg496 <= $signed({{$unsigned({reg457, reg458}), reg485},
              $signed($unsigned(reg458[(1'h0):(1'h0)]))});
          if ($unsigned((8'hb3)))
            begin
              reg497 <= $signed((reg493[(4'h9):(4'h8)] ^ $unsigned(reg477)));
              reg498 <= reg451;
              reg499 = $signed($signed((!reg469[(5'h10):(4'h9)])));
              reg500 = reg497[(2'h2):(2'h2)];
            end
          else
            begin
              reg499 = $signed(reg442);
              reg501 <= wire435;
              reg502 = $unsigned(((~&$unsigned({reg437})) ?
                  $unsigned(reg496) : reg458));
            end
          for (forvar503 = (1'h0); (forvar503 < (2'h2)); forvar503 = (forvar503 + (1'h1)))
            begin
              reg504 = {$unsigned(((~^(~|reg469)) << $unsigned(wire433[(4'hf):(4'h9)])))};
              reg505 = (&reg486[(1'h0):(1'h0)]);
              reg506 <= reg450[(1'h1):(1'h1)];
              reg507 = (reg474 ?
                  $unsigned(reg481) : (reg495 ?
                      $signed({$signed(reg461),
                          reg440}) : $unsigned({reg504[(4'ha):(4'h8)]})));
            end
          reg508 <= (-(reg446 ?
              (7'h4a) : (+((-wire464) ?
                  $unsigned(reg488) : (reg446 ? wire435 : reg506)))));
        end
      else
        begin
          if ((8'ha4))
            begin
              reg499 = forvar503[(2'h2):(2'h2)];
              reg501 <= ((reg437[(3'h4):(1'h1)] ^~ $signed(((reg461 | reg446) > reg459))) ?
                  ((((^~reg440) < (wire464 * reg486)) ^~ reg497) ?
                      reg486 : reg439[(4'h9):(3'h6)]) : reg481);
              reg503 <= {reg485[(4'h9):(4'h8)]};
              reg504 = (~^({(&$unsigned((8'ha6)))} ?
                  (({reg485} ? (~&reg494) : (reg481 ? reg451 : reg496)) ?
                      $unsigned(reg494[(4'hb):(1'h0)]) : (reg451 ?
                          (reg458 <<< reg503) : reg504[(3'h7):(1'h1)])) : reg508));
            end
          else
            begin
              reg495 <= ($unsigned({(-$unsigned(reg490)),
                  $unsigned($unsigned(wire465))}) >= wire429[(2'h3):(1'h1)]);
            end
          for (forvar505 = (1'h0); (forvar505 < (1'h0)); forvar505 = (forvar505 + (1'h1)))
            begin
              reg506 <= (wire434 ?
                  reg494[(5'h15):(4'he)] : (((~|reg505) ?
                      reg497 : $signed((forvar503 ?
                          wire464 : reg503))) >> (-(+$signed(reg494)))));
              reg507 = ({reg439[(5'h13):(1'h1)]} ?
                  (((reg502[(2'h3):(1'h0)] < (8'ha2)) & (reg471[(4'ha):(4'h8)] > (~&reg504))) <= $unsigned(((~&reg471) ?
                      (^~reg494) : (reg486 ^~ reg506)))) : forvar503);
              reg509 = (8'hb9);
            end
          reg510 <= $unsigned(($signed(((8'ha2) ?
                  wire435[(3'h4):(2'h2)] : reg499)) ?
              forvar503 : reg505[(1'h0):(1'h0)]));
          for (forvar511 = (1'h0); (forvar511 < (1'h1)); forvar511 = (forvar511 + (1'h1)))
            begin
              reg512 <= $signed((reg442[(3'h7):(3'h6)] ?
                  {{wire435[(3'h4):(1'h0)],
                          reg504}} : $signed($signed((wire429 ?
                      reg499 : wire464)))));
              reg513 = (+(reg498[(5'h10):(1'h0)] ?
                  reg442[(4'ha):(2'h3)] : $signed($unsigned((wire435 ?
                      reg496 : reg508)))));
              reg514 = $signed($signed($unsigned(reg485)));
              reg515 = (($signed($signed(reg497[(2'h3):(1'h0)])) >> $unsigned(($signed(reg512) < (reg499 ?
                  wire464 : reg490)))) != reg485);
              reg516 = $signed(($unsigned($unsigned((&reg514))) ?
                  ((-$signed(wire435)) ^ reg477[(4'h9):(3'h4)]) : {reg485,
                      (reg502 & reg503[(3'h7):(3'h5)])}));
            end
          reg517 = wire432;
        end
      if (((reg506 ^ reg514[(1'h1):(1'h1)]) + (~^reg496[(4'hb):(3'h5)])))
        begin
          reg518 <= {(~wire429[(2'h2):(1'h0)])};
          for (forvar519 = (1'h0); (forvar519 < (1'h0)); forvar519 = (forvar519 + (1'h1)))
            begin
              reg520 <= wire433[(4'he):(4'h9)];
              reg521 = $unsigned(reg493[(2'h3):(2'h3)]);
              reg522 = (!(~|{(((8'ha5) ?
                      reg513 : reg514) && reg500[(4'h9):(2'h3)])}));
            end
          if ($signed($unsigned($unsigned({$signed((8'haf)),
              $signed(reg503)}))))
            begin
              reg523 = (($signed(reg505) || $unsigned($signed(reg438[(1'h1):(1'h0)]))) ^~ (8'ha4));
              reg524 = (8'hb4);
              reg525 <= (forvar519 >= {$unsigned((-$unsigned((7'h46)))),
                  {(reg515 ? reg516[(1'h1):(1'h1)] : ((8'h9f) >= reg488))}});
            end
          else
            begin
              reg525 <= {$unsigned({$signed((~&reg488))}), $unsigned((7'h47))};
              reg526 <= $signed({reg458[(2'h3):(2'h2)],
                  (($unsigned(reg486) > (-reg451)) + forvar519[(2'h3):(2'h3)])});
              reg527 <= ($unsigned($signed($unsigned((reg525 ?
                      reg488 : reg491)))) ?
                  ($signed((wire430 ?
                      (wire432 ?
                          reg437 : reg510) : (forvar503 <<< reg439))) ^~ (wire465[(5'h14):(3'h4)] && ((wire433 ^ wire434) - reg490[(5'h18):(5'h14)]))) : $signed(reg450));
              reg528 <= reg496[(4'he):(4'hb)];
              reg529 <= reg498[(3'h4):(3'h4)];
            end
          if ((forvar503[(1'h0):(1'h0)] != ((8'hbc) ?
              (^(|((8'hae) ?
                  reg439 : reg517))) : $signed(((wire434 != forvar505) ?
                  ((7'h4a) ? reg491 : reg527) : $signed(reg507))))))
            begin
              reg530 = wire431;
              reg531 <= wire464;
              reg532 <= (^$signed($unsigned(($signed(reg459) + reg527[(1'h0):(1'h0)]))));
              reg533 <= (reg523[(1'h0):(1'h0)] ?
                  wire465 : (reg438 ?
                      reg522[(1'h1):(1'h0)] : ($signed(reg515[(4'hb):(1'h1)]) ?
                          $signed($unsigned(reg491)) : $unsigned(reg509))));
            end
          else
            begin
              reg531 <= reg496;
              reg534 = reg486;
              reg535 = $signed(((+$unsigned((8'ha5))) ?
                  ((reg523 || ((7'h47) - reg507)) ?
                      (((8'hb3) * reg495) ~^ (reg494 == forvar511)) : reg502) : wire435[(1'h1):(1'h1)]));
            end
        end
      else
        begin
          for (forvar518 = (1'h0); (forvar518 < (2'h3)); forvar518 = (forvar518 + (1'h1)))
            begin
              reg519 <= (&(wire431 ?
                  $unsigned($signed($unsigned(reg535))) : {{$unsigned((8'hb0)),
                          $unsigned(reg494)}}));
              reg520 <= $unsigned($signed(reg488[(2'h3):(1'h1)]));
              reg525 <= (reg529[(1'h1):(1'h0)] ?
                  (((7'h4a) ?
                      ((~&reg526) + $unsigned(reg500)) : $signed($signed(reg517))) ^ $unsigned({$signed(reg477),
                      $unsigned(reg531)})) : reg503);
            end
          for (forvar526 = (1'h0); (forvar526 < (2'h2)); forvar526 = (forvar526 + (1'h1)))
            begin
              reg530 = $unsigned(wire464);
              reg531 <= $signed(reg507[(3'h4):(3'h4)]);
              reg532 <= reg439[(2'h3):(1'h1)];
            end
          reg533 <= reg481[(3'h7):(3'h6)];
        end
      for (forvar536 = (1'h0); (forvar536 < (2'h2)); forvar536 = (forvar536 + (1'h1)))
        begin
          reg537 = $unsigned($signed((reg521 ~^ {$signed(wire432)})));
          if (reg440)
            begin
              reg538 = {(reg507[(1'h0):(1'h0)] <= ((&reg529[(4'hb):(1'h1)]) * ((8'ha3) ?
                      (!wire431) : reg493)))};
              reg539 = ($unsigned(reg481[(2'h2):(2'h2)]) | forvar505[(4'he):(1'h1)]);
              reg540 <= $signed(forvar519[(4'hc):(2'h3)]);
              reg541 = {(wire465[(5'h12):(3'h7)] ?
                      reg539[(4'h8):(1'h1)] : $unsigned($signed($unsigned(wire435)))),
                  {{($signed(reg515) ? (8'h9c) : ((8'haf) ? reg469 : (8'ha3))),
                          reg527[(3'h5):(3'h5)]}}};
              reg542 <= (($unsigned(reg477) ?
                  $signed((reg451[(3'h5):(1'h0)] ?
                      reg512 : (~|reg510))) : reg461[(4'h8):(4'h8)]) < (^~reg524[(5'h17):(3'h5)]));
            end
          else
            begin
              reg540 <= $signed($unsigned(((forvar519 >>> reg540) || reg442)));
              reg542 <= ((reg491[(3'h4):(2'h2)] ?
                  ((reg512 != (reg535 >>> reg531)) & (+wire429[(2'h2):(1'h1)])) : $signed((~reg508[(3'h6):(2'h3)]))) + reg519[(2'h3):(1'h1)]);
              reg543 = reg469[(4'h8):(2'h2)];
              reg544 <= $unsigned((wire434[(3'h5):(2'h2)] ?
                  reg494 : $signed(reg450[(1'h0):(1'h0)])));
            end
          for (forvar545 = (1'h0); (forvar545 < (3'h4)); forvar545 = (forvar545 + (1'h1)))
            begin
              reg546 = (reg491[(2'h3):(1'h1)] <<< $signed((~$unsigned((|(7'h48))))));
              reg547 <= (^~$signed((reg437[(2'h2):(1'h0)] > $unsigned(reg512))));
              reg548 = reg494[(4'hb):(3'h6)];
              reg549 <= {(8'hb5)};
            end
        end
      for (forvar550 = (1'h0); (forvar550 < (3'h4)); forvar550 = (forvar550 + (1'h1)))
        begin
          for (forvar551 = (1'h0); (forvar551 < (2'h3)); forvar551 = (forvar551 + (1'h1)))
            begin
              reg552 <= $signed((~$unsigned((|$signed(wire465)))));
              reg553 <= $signed((~^(((^~reg494) ^~ {reg442}) ?
                  (reg498 > (reg496 ? reg491 : reg541)) : reg481)));
              reg554 = (((8'ha5) ?
                      (reg509 ?
                          (~|(reg439 - forvar526)) : ($unsigned(reg543) ?
                              forvar503[(1'h1):(1'h0)] : forvar519[(1'h1):(1'h1)])) : $unsigned(forvar505[(4'hf):(1'h0)])) ?
                  (($unsigned(((7'h40) ? reg552 : (8'hbd))) ?
                          (!forvar551[(2'h2):(1'h0)]) : reg469) ?
                      $signed($signed((reg459 ?
                          reg539 : reg524))) : ($unsigned(reg481[(2'h2):(2'h2)]) ?
                          {(|reg553)} : reg534)) : (reg529 ?
                      reg504[(4'h9):(3'h4)] : reg530[(3'h4):(2'h2)]));
              reg555 <= reg527[(3'h6):(3'h6)];
            end
          if ($signed((reg527 << (8'hb0))))
            begin
              reg556 = ({({forvar550[(1'h1):(1'h0)]} ?
                          reg529[(3'h6):(1'h1)] : forvar518[(3'h6):(3'h6)]),
                      $signed($unsigned((!reg518)))} ?
                  $signed($signed($signed($unsigned(reg520)))) : (forvar511 ?
                      $unsigned(reg508) : (&$signed((^~reg518)))));
              reg557 <= $signed(((({reg498,
                  reg471} >>> forvar518) <= $signed((|forvar545))) >>> (reg520 ?
                  {wire430, reg510} : (+(!reg526)))));
            end
          else
            begin
              reg556 = (reg515 << {$signed((~|{reg525, (8'hbf)})),
                  (|(((8'hb3) ? reg537 : reg461) ?
                      forvar526[(2'h2):(1'h1)] : $signed(reg513)))});
              reg558 = reg469[(5'h15):(4'h8)];
              reg559 = (($signed((~|((8'hb5) * (8'ha1)))) * ($unsigned((|reg529)) || $signed({forvar551,
                      reg552}))) ?
                  {$unsigned(((-(8'h9e)) ?
                          (reg516 < (8'hb1)) : $unsigned((8'h9d)))),
                      wire432[(1'h1):(1'h0)]} : ((reg513[(1'h1):(1'h1)] != (~&(reg546 ?
                          (8'ha5) : reg553))) ?
                      ((8'hbc) ?
                          $signed((8'hb3)) : (reg523[(1'h0):(1'h0)] != reg437[(1'h1):(1'h0)])) : $unsigned((~&(^(7'h4a))))));
              reg560 <= wire433[(4'h9):(1'h1)];
              reg561 = reg496;
            end
          for (forvar562 = (1'h0); (forvar562 < (3'h4)); forvar562 = (forvar562 + (1'h1)))
            begin
              reg563 <= (^~reg438[(3'h7):(1'h0)]);
            end
          reg564 = reg500;
        end
      reg565 = $unsigned($signed((^($signed(forvar519) ?
          (reg438 ? (8'hb8) : reg546) : reg437))));
    end
  assign wire566 = $signed(reg494);
  assign wire567 = $signed(reg469);
  always
    @(posedge clk) begin
      for (forvar568 = (1'h0); (forvar568 < (1'h0)); forvar568 = (forvar568 + (1'h1)))
        begin
          for (forvar569 = (1'h0); (forvar569 < (1'h1)); forvar569 = (forvar569 + (1'h1)))
            begin
              reg570 = {reg442};
            end
          reg571 <= wire432;
          if (($unsigned($unsigned(((reg490 ^~ (7'h45)) ^ (reg474 * reg442)))) >> (+{$unsigned($unsigned(reg552))})))
            begin
              reg572 = reg469[(4'ha):(3'h6)];
              reg573 = $signed(reg495[(3'h6):(3'h4)]);
              reg574 = $signed(((7'h4a) ?
                  $unsigned(($unsigned(reg529) ?
                      reg438 : $unsigned(wire465))) : $unsigned(($unsigned(reg495) <<< reg498[(3'h6):(2'h2)]))));
            end
          else
            begin
              reg575 <= reg498;
              reg576 = {$unsigned((($unsigned(reg575) < reg575) + $signed(reg508)))};
              reg577 = $unsigned(($unsigned(reg491) && (8'hb7)));
              reg578 <= $unsigned($unsigned((~|$signed($signed((7'h43))))));
              reg579 = wire465;
            end
        end
      if (((^~($signed((~&reg533)) ?
              $unsigned($unsigned(reg560)) : $unsigned($unsigned(reg503)))) ?
          reg481 : (^~$signed($unsigned($unsigned(reg572))))))
        begin
          for (forvar580 = (1'h0); (forvar580 < (2'h3)); forvar580 = (forvar580 + (1'h1)))
            begin
              reg581 = reg532;
              reg582 <= reg494[(5'h14):(4'h9)];
              reg583 = ($unsigned((&reg557[(2'h3):(1'h1)])) ?
                  ({((8'haa) > $signed(reg575)),
                          ($unsigned(reg529) ? $signed(reg490) : reg519)} ?
                      $signed((~^$signed(reg582))) : (reg576[(5'h10):(4'hd)] || reg490[(2'h3):(2'h2)])) : (~$unsigned(reg547[(2'h3):(2'h3)])));
              reg584 <= $signed((({(~reg459)} ?
                  {reg450[(1'h0):(1'h0)], {(8'ha7), reg542}} : ((reg583 ?
                      reg571 : wire465) || (reg540 ?
                      reg493 : reg469))) == reg525[(4'h8):(3'h5)]));
            end
          if (($unsigned(reg572) ?
              $signed((((~reg485) << (8'ha0)) ?
                  (reg532[(4'he):(3'h7)] && $signed(reg446)) : ((8'haa) ?
                      $signed((8'ha8)) : $signed(reg494)))) : reg488[(3'h6):(1'h1)]))
            begin
              reg585 = (+$unsigned($unsigned($signed((reg581 * reg457)))));
            end
          else
            begin
              reg586 <= ({reg572} ?
                  $signed((+((wire431 ? reg526 : wire431) ?
                      (reg519 ?
                          reg442 : reg572) : reg477))) : {$unsigned({reg542})});
              reg587 = reg442[(2'h3):(1'h0)];
              reg588 <= $signed($signed(reg506));
              reg589 <= (reg560 ?
                  $unsigned((((reg490 <<< wire434) >>> {reg553}) > (|$unsigned(reg498)))) : (^~reg572[(3'h7):(3'h7)]));
              reg590 = $signed(reg586);
            end
          reg591 = reg481;
          if ((($signed(reg573) ^~ (8'hbf)) == {reg528[(4'ha):(4'ha)]}))
            begin
              reg592 <= ((($signed(((8'ha9) ?
                          reg510 : reg540)) <<< ($unsigned(reg510) ?
                          {(7'h48), reg532} : $signed((8'hb5)))) ?
                      (8'hbb) : (reg540[(4'hb):(2'h2)] ?
                          (^reg542) : $signed($signed(reg446)))) ?
                  reg518 : $unsigned({{(reg581 ? (8'hb1) : reg553), reg540},
                      $unsigned((wire566 ? reg549 : reg552))}));
              reg593 = {$unsigned((!(^reg503))),
                  ((((reg494 > reg575) | {reg493, reg510}) <= reg451) ?
                      $unsigned($unsigned($unsigned(reg579))) : $signed(((reg506 ?
                          wire430 : reg529) == $unsigned(reg549))))};
            end
          else
            begin
              reg592 <= reg533[(3'h5):(2'h3)];
              reg593 = ((((~&(reg590 ? reg588 : (8'hbe))) ?
                          reg488[(2'h3):(1'h1)] : $unsigned({reg501})) ?
                      $signed($signed(((8'had) + reg573))) : reg493[(1'h0):(1'h0)]) ?
                  (~($unsigned(reg459) ?
                      (reg573[(4'h9):(3'h4)] ?
                          reg519[(2'h3):(1'h1)] : reg584) : reg533)) : reg437[(3'h4):(2'h2)]);
              reg594 <= $signed(($unsigned($unsigned(reg481)) ?
                  $signed((reg440 ?
                      reg573 : $unsigned(reg461))) : $unsigned(reg590[(3'h7):(1'h1)])));
              reg595 = reg552;
            end
          if ((wire464 || {reg570[(1'h0):(1'h0)]}))
            begin
              reg596 = $unsigned($unsigned((reg520[(1'h0):(1'h0)] ?
                  reg459 : (^$unsigned(reg520)))));
              reg597 = (^$signed($signed($unsigned($unsigned(reg520)))));
              reg598 = reg542;
              reg599 <= ($unsigned((reg510[(2'h3):(1'h1)] ?
                      wire429[(3'h4):(1'h0)] : ((8'hae) || $signed(reg527)))) ?
                  reg471 : $signed(($signed((+wire433)) ?
                      reg497[(2'h2):(1'h0)] : reg529[(2'h3):(1'h1)])));
              reg600 <= (reg526[(4'h9):(3'h6)] < $unsigned((-$signed(reg525[(4'h8):(4'h8)]))));
            end
          else
            begin
              reg599 <= (reg557 ?
                  (reg496[(4'hd):(3'h7)] ?
                      $signed(wire465[(4'hc):(3'h4)]) : $signed($signed(wire430))) : ((reg576[(4'h8):(3'h6)] ?
                      (-(reg549 ~^ reg451)) : wire433[(3'h5):(1'h0)]) + ({(reg581 || (8'hba)),
                      ((7'h49) >= reg493)} + ({(8'had),
                      (8'haf)} || (~(8'hab))))));
              reg601 = ((~((8'hae) ^~ reg519)) ?
                  $unsigned((^~$signed($signed(wire465)))) : ((!reg575[(3'h7):(3'h6)]) >= $unsigned($unsigned($unsigned(reg481)))));
              reg602 = (+$signed($signed($unsigned($signed(reg486)))));
            end
        end
      else
        begin
          for (forvar580 = (1'h0); (forvar580 < (1'h1)); forvar580 = (forvar580 + (1'h1)))
            begin
              reg582 <= $signed(($unsigned(reg591) <<< (7'h4a)));
              reg583 = $signed(($signed((&(|reg510))) ?
                  (reg508 ?
                      reg485 : ((~|reg491) <= (!reg528))) : ($unsigned((~&reg596)) > reg542)));
              reg584 <= reg474;
            end
        end
      reg603 <= ((&(!($signed(wire465) ?
          reg474[(4'ha):(3'h6)] : (|reg531)))) >>> $signed((($unsigned(wire464) == wire432[(3'h6):(1'h0)]) < (^(reg601 >> reg508)))));
      if ((((+reg440[(2'h2):(1'h0)]) > (~|((^forvar568) ?
          (^reg481) : reg496))) && $signed((reg560[(4'hc):(4'hc)] ?
          wire430 : ($signed(reg508) <<< $signed(reg595))))))
        begin
          if ($signed($unsigned(reg533)))
            begin
              reg604 <= (~&reg519);
              reg605 = $unsigned({(($signed(reg495) <<< reg457[(2'h2):(1'h1)]) != (|(reg477 ?
                      reg599 : wire566)))});
              reg606 = wire435[(2'h3):(2'h2)];
              reg607 <= reg439[(5'h12):(2'h2)];
              reg608 <= (({reg587,
                      (reg528[(3'h6):(3'h6)] ?
                          reg532 : reg490[(4'he):(3'h7)])} ?
                  reg503[(5'h13):(4'ha)] : (8'hbc)) != ((reg540 << $unsigned((reg457 ?
                  reg450 : (8'hab)))) & $signed(({(8'hbe),
                  reg512} >= $unsigned(reg557)))));
            end
          else
            begin
              reg604 <= $unsigned((reg557[(4'h8):(3'h4)] | $unsigned((reg442[(2'h2):(1'h1)] ^ (reg437 - reg557)))));
              reg607 <= reg496[(3'h4):(2'h2)];
              reg608 <= $unsigned((-reg601));
              reg609 = ((({(reg440 ?
                              reg457 : wire464)} >> reg469[(3'h6):(1'h0)]) ?
                      reg589 : reg582) ?
                  (wire433 ?
                      (+$signed(wire433[(1'h1):(1'h1)])) : reg495) : (8'hbd));
              reg610 <= $signed($unsigned(reg494));
            end
          reg611 <= reg589;
          if (reg582[(2'h3):(2'h2)])
            begin
              reg612 <= ($signed(reg498) ?
                  reg555[(3'h5):(1'h0)] : (!($unsigned($unsigned(reg555)) <= $signed((reg497 <<< reg563)))));
              reg613 <= reg608[(2'h2):(1'h1)];
              reg614 = reg544[(3'h4):(2'h2)];
              reg615 = {reg526[(4'ha):(2'h3)], reg608[(2'h2):(1'h0)]};
              reg616 = reg519;
            end
          else
            begin
              reg614 = $signed(((reg437[(2'h3):(1'h0)] ?
                  reg450 : reg574[(2'h2):(1'h0)]) ^ (-(!(|wire567)))));
              reg615 = $signed(reg579[(5'h10):(3'h4)]);
              reg616 = $signed($unsigned(reg525));
              reg617 = reg442;
              reg618 = ((reg560[(4'ha):(2'h2)] >= reg575[(3'h4):(2'h2)]) ?
                  $unsigned($signed(($unsigned(reg528) ?
                      ((8'hbd) - reg615) : (reg585 ?
                          reg607 : reg603)))) : $unsigned(reg533));
            end
        end
      else
        begin
          reg604 <= reg442;
          reg607 <= reg490[(1'h1):(1'h0)];
          if ($unsigned((&(reg485 > (reg615 ? $unsigned(reg605) : reg529)))))
            begin
              reg609 = reg477;
              reg610 <= $signed(((8'ha2) ?
                  reg597[(3'h5):(1'h0)] : (+{(~(8'ha2))})));
              reg611 <= (reg540 ^~ ($signed(reg494) - (8'hac)));
              reg614 = (reg533 ?
                  (((8'ha2) ^~ $unsigned((reg603 > reg503))) ^~ $unsigned($signed((reg450 + (8'hb6))))) : reg588[(4'h9):(2'h2)]);
              reg615 = $unsigned($signed($unsigned((&(reg577 ?
                  wire465 : reg469)))));
            end
          else
            begin
              reg608 <= $unsigned({($signed($signed((8'hbb))) > reg611[(4'hd):(4'h8)])});
              reg609 = $signed(reg461[(5'h11):(3'h6)]);
              reg614 = ($signed($signed(reg618)) ?
                  (-$unsigned((8'hbf))) : wire465[(4'hf):(1'h1)]);
              reg619 <= reg584;
              reg620 <= $unsigned((^~(|reg438[(4'h9):(3'h7)])));
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module394  (y, clk, wire398, wire397, wire396, wire395);
  output wire [(32'h172):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire398;
  input wire [(5'h13):(1'h0)] wire397;
  input wire signed [(3'h5):(1'h0)] wire396;
  input wire [(3'h6):(1'h0)] wire395;
  wire [(4'hc):(1'h0)] wire425;
  wire [(5'h10):(1'h0)] wire424;
  wire signed [(4'h9):(1'h0)] wire399;
  reg [(5'h10):(1'h0)] reg423 = (1'h0);
  reg [(5'h18):(1'h0)] reg414 = (1'h0);
  reg [(3'h4):(1'h0)] reg411 = (1'h0);
  reg [(2'h3):(1'h0)] reg410 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg407 = (1'h0);
  reg [(5'h17):(1'h0)] reg406 = (1'h0);
  reg [(4'ha):(1'h0)] reg405 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg401 = (1'h0);
  reg [(5'h17):(1'h0)] reg400 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg422 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg421 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg420 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg419 = (1'h0);
  reg signed [(4'he):(1'h0)] reg418 = (1'h0);
  reg [(5'h12):(1'h0)] reg417 = (1'h0);
  reg [(4'hb):(1'h0)] reg416 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg415 = (1'h0);
  reg [(5'h11):(1'h0)] forvar413 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg412 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg409 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar408 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg404 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg403 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg402 = (1'h0);
  assign y = {wire425,
                 wire424,
                 wire399,
                 reg423,
                 reg414,
                 reg411,
                 reg410,
                 reg407,
                 reg406,
                 reg405,
                 reg401,
                 reg400,
                 reg422,
                 reg421,
                 reg420,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 forvar413,
                 reg412,
                 reg409,
                 forvar408,
                 reg404,
                 reg403,
                 reg402,
                 (1'h0)};
  assign wire399 = $unsigned($signed(((^~wire396[(2'h3):(2'h3)]) << ($signed((8'ha3)) == wire397))));
  always
    @(posedge clk) begin
      reg400 <= $unsigned({(wire399[(4'h9):(1'h1)] ?
              $signed(wire395) : ($signed(wire395) ?
                  (wire398 ? (8'hac) : wire395) : (wire399 ?
                      wire395 : wire397)))});
      if ($unsigned({$unsigned(wire398[(3'h6):(2'h2)])}))
        begin
          if ((|wire397[(4'ha):(3'h5)]))
            begin
              reg401 <= (({(((8'hbb) ? reg400 : wire397) == (wire395 ?
                          (8'hab) : reg400))} ?
                  wire397[(4'hd):(1'h1)] : ((wire399[(2'h2):(1'h1)] ?
                          reg400 : $signed((7'h47))) ?
                      {(~^reg400)} : ((|wire396) ^~ reg400[(1'h0):(1'h0)]))) + wire397);
            end
          else
            begin
              reg401 <= (wire396 ?
                  {$unsigned(((reg401 ?
                          wire395 : reg400) - $unsigned((7'h40)))),
                      reg400[(3'h5):(2'h3)]} : $signed(wire396[(2'h3):(1'h0)]));
            end
          reg402 = $unsigned(((wire399 ?
                  (wire398 ?
                      (~&wire399) : $unsigned(wire395)) : $unsigned((+wire398))) ?
              (($signed(wire397) ? (!wire399) : (wire395 ? reg400 : wire398)) ?
                  wire396 : ({wire399, reg401} ?
                      {wire398} : (reg400 ? wire397 : reg400))) : {((wire395 ?
                      reg400 : wire397) > (reg400 ? wire399 : reg401))}));
          reg403 = reg401;
          reg404 = $signed($signed(($signed(wire396[(1'h1):(1'h1)]) ?
              (wire399[(1'h1):(1'h1)] * (reg402 ?
                  wire399 : wire399)) : (&$unsigned(reg400)))));
        end
      else
        begin
          if ($unsigned($unsigned(((+(^~reg404)) | (8'ha5)))))
            begin
              reg401 <= reg401[(4'hb):(1'h0)];
              reg405 <= $signed(reg404[(2'h3):(1'h1)]);
            end
          else
            begin
              reg402 = ($unsigned($signed({{reg405, wire397}})) ?
                  $signed((~|((^(8'hb3)) ?
                      (wire396 ?
                          wire399 : reg402) : reg402[(2'h2):(2'h2)]))) : ((wire397 + ({wire396,
                              reg402} ?
                          $unsigned(wire399) : (wire396 >> (8'ha1)))) ?
                      $signed(($unsigned(reg405) ~^ (reg403 ?
                          reg401 : reg403))) : $unsigned(reg400[(2'h3):(2'h2)])));
              reg403 = $signed((8'haa));
              reg405 <= (wire397 ?
                  reg402 : $signed((^~((wire399 ?
                      (8'hb4) : (7'h48)) + $unsigned(reg401)))));
              reg406 <= reg400;
              reg407 <= (($unsigned(reg406) ?
                      (~^$signed(reg404[(2'h2):(2'h2)])) : $unsigned({(reg402 ?
                              reg401 : (8'ha5)),
                          $unsigned(reg405)})) ?
                  $signed((reg404 ^ $signed(((7'h40) ?
                      wire396 : reg402)))) : (|(wire397[(4'he):(2'h3)] + wire399[(3'h5):(3'h5)])));
            end
          for (forvar408 = (1'h0); (forvar408 < (2'h2)); forvar408 = (forvar408 + (1'h1)))
            begin
              reg409 = (-(!(($unsigned(wire395) ?
                  $unsigned(wire398) : $signed(wire395)) ^~ wire399)));
              reg410 <= (((($unsigned(reg406) ?
                      reg401[(4'h9):(2'h3)] : {(7'h47), wire396}) < (|reg404)) ?
                  wire398 : (~$signed({reg405,
                      forvar408}))) || $signed(($unsigned(wire399) | ((reg403 ?
                  reg405 : forvar408) + (wire398 << reg409)))));
            end
          reg411 <= (($signed($unsigned($unsigned(reg407))) ?
                  (!(^~(7'h46))) : $unsigned(reg410)) ?
              reg407[(4'ha):(3'h7)] : (~{((+forvar408) ?
                      $signed(reg403) : $unsigned((8'hbd)))}));
          reg412 = $signed(reg405);
          for (forvar413 = (1'h0); (forvar413 < (3'h4)); forvar413 = (forvar413 + (1'h1)))
            begin
              reg414 <= ({wire399[(4'h8):(4'h8)]} && {$signed(reg411)});
              reg415 = ((^reg414[(4'hb):(2'h3)]) != ((reg407[(4'hf):(4'hf)] ?
                  $unsigned((8'hab)) : ($signed(reg411) ?
                      $unsigned(reg405) : (~reg406))) << reg410[(2'h3):(2'h2)]));
              reg416 = (^reg414);
              reg417 = (~&$signed((8'ha3)));
              reg418 = ((reg401 ?
                  ($unsigned($unsigned(reg402)) ?
                      ($signed(reg403) ?
                          reg404[(5'h12):(1'h0)] : $signed(wire397)) : reg416[(3'h7):(3'h7)]) : ({reg405[(3'h6):(3'h6)],
                      $signed(reg406)} ~^ ((~&reg415) ?
                      $signed((8'ha5)) : $signed(reg409)))) != {(~^(reg402 ?
                      reg409[(4'hc):(3'h6)] : $signed(reg411))),
                  (^$signed(((8'ha3) ? reg407 : (7'h40))))});
            end
        end
    end
  always
    @(posedge clk) begin
      reg419 = (reg410[(1'h1):(1'h0)] >>> ($unsigned(($signed(wire396) >> wire397)) ?
          reg410[(2'h3):(2'h2)] : $signed({$signed((7'h41)), (~&reg414)})));
      reg420 = (($unsigned(((wire395 << reg411) ?
          reg401 : (reg414 ^ wire398))) & $signed(($unsigned(reg411) ?
          reg401 : (~|reg405)))) << ((~&reg401) * $unsigned($signed((-reg406)))));
      reg421 = reg407;
      reg422 = (reg420 ?
          wire395[(1'h0):(1'h0)] : (($unsigned((~^reg405)) ?
                  reg407 : ((~|reg406) ? (8'hb1) : reg400)) ?
              ($signed((|reg420)) != $unsigned((reg421 ?
                  reg400 : reg407))) : ((8'h9e) ?
                  $unsigned($signed((8'hbc))) : (8'hb0))));
      reg423 <= wire397[(4'hf):(4'h9)];
    end
  assign wire424 = (($signed((8'ha6)) * {(~|(!wire398))}) ?
                       wire398 : (~({$unsigned(wire397)} ?
                           reg401[(1'h1):(1'h1)] : reg423)));
  assign wire425 = (-{reg405, $signed({$unsigned((8'hbd))})});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1192
#(parameter param1287 = ((((^~(8'hac)) && (~((8'haa) || (8'hb1)))) ? (7'h42) : ((~(~|(8'hb1))) ? ((-(8'ha3)) ? ((8'hae) >>> (8'hac)) : (8'hbb)) : ((&(8'hbb)) && (^~(7'h48))))) << (((&((7'h45) ? (8'ha8) : (8'hb6))) >>> {{(7'h48)}}) < (({(7'h44)} ? {(8'haf)} : (~&(8'hbd))) ? ({(7'h47), (8'hbf)} < ((8'h9c) ? (7'h40) : (8'hb8))) : (8'hab)))))
(y, clk, wire1197, wire1196, wire1195, wire1194, wire1193);
  output wire [(32'h4b4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h15):(1'h0)] wire1197;
  input wire signed [(4'he):(1'h0)] wire1196;
  input wire [(5'h13):(1'h0)] wire1195;
  input wire signed [(5'h16):(1'h0)] wire1194;
  input wire signed [(5'h13):(1'h0)] wire1193;
  wire [(4'h8):(1'h0)] wire1212;
  wire signed [(5'h15):(1'h0)] wire1211;
  reg [(5'h12):(1'h0)] reg1284 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1283 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1282 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1280 = (1'h0);
  reg [(4'ha):(1'h0)] reg1278 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1276 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1266 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1265 = (1'h0);
  reg [(4'he):(1'h0)] reg1263 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1258 = (1'h0);
  reg [(4'hb):(1'h0)] reg1257 = (1'h0);
  reg [(5'h17):(1'h0)] reg1254 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1253 = (1'h0);
  reg [(5'h18):(1'h0)] reg1251 = (1'h0);
  reg [(5'h14):(1'h0)] reg1250 = (1'h0);
  reg [(4'he):(1'h0)] reg1249 = (1'h0);
  reg [(4'h9):(1'h0)] reg1248 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1246 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1245 = (1'h0);
  reg [(3'h6):(1'h0)] reg1243 = (1'h0);
  reg [(4'ha):(1'h0)] reg1238 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1235 = (1'h0);
  reg [(5'h13):(1'h0)] reg1230 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1229 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1226 = (1'h0);
  reg [(2'h3):(1'h0)] reg1223 = (1'h0);
  reg [(5'h14):(1'h0)] reg1222 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1219 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1218 = (1'h0);
  reg [(4'h8):(1'h0)] reg1217 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1214 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1213 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1210 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1209 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1207 = (1'h0);
  reg [(5'h13):(1'h0)] reg1205 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1204 = (1'h0);
  reg [(4'h9):(1'h0)] reg1199 = (1'h0);
  reg [(2'h3):(1'h0)] reg1200 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1286 = (1'h0);
  reg [(3'h4):(1'h0)] reg1285 = (1'h0);
  reg [(2'h2):(1'h0)] reg1281 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1279 = (1'h0);
  reg [(5'h17):(1'h0)] reg1277 = (1'h0);
  reg [(5'h12):(1'h0)] reg1275 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1274 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1273 = (1'h0);
  reg [(4'he):(1'h0)] reg1272 = (1'h0);
  reg [(4'he):(1'h0)] reg1271 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1270 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1269 = (1'h0);
  reg [(3'h5):(1'h0)] reg1268 = (1'h0);
  reg [(2'h3):(1'h0)] reg1267 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1264 = (1'h0);
  reg [(3'h4):(1'h0)] reg1262 = (1'h0);
  reg [(5'h18):(1'h0)] reg1261 = (1'h0);
  reg [(5'h14):(1'h0)] reg1260 = (1'h0);
  reg [(3'h7):(1'h0)] reg1259 = (1'h0);
  reg [(4'ha):(1'h0)] reg1256 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1255 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1252 = (1'h0);
  reg [(4'ha):(1'h0)] reg1247 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1244 = (1'h0);
  reg [(5'h13):(1'h0)] reg1242 = (1'h0);
  reg [(5'h16):(1'h0)] reg1241 = (1'h0);
  reg [(3'h7):(1'h0)] reg1240 = (1'h0);
  reg [(4'h8):(1'h0)] reg1239 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1237 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1236 = (1'h0);
  reg [(5'h16):(1'h0)] reg1234 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1233 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar1232 = (1'h0);
  reg [(5'h15):(1'h0)] reg1231 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1228 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1227 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1225 = (1'h0);
  reg [(2'h2):(1'h0)] reg1224 = (1'h0);
  reg [(5'h13):(1'h0)] forvar1221 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1220 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1216 = (1'h0);
  reg [(3'h4):(1'h0)] reg1215 = (1'h0);
  reg [(5'h15):(1'h0)] reg1208 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1206 = (1'h0);
  reg [(5'h14):(1'h0)] reg1203 = (1'h0);
  reg [(5'h15):(1'h0)] reg1202 = (1'h0);
  reg [(5'h12):(1'h0)] reg1201 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1199 = (1'h0);
  reg [(5'h13):(1'h0)] reg1198 = (1'h0);
  assign y = {wire1212,
                 wire1211,
                 reg1284,
                 reg1283,
                 reg1282,
                 reg1280,
                 reg1278,
                 reg1276,
                 reg1266,
                 reg1265,
                 reg1263,
                 reg1258,
                 reg1257,
                 reg1254,
                 reg1253,
                 reg1251,
                 reg1250,
                 reg1249,
                 reg1248,
                 reg1246,
                 reg1245,
                 reg1243,
                 reg1238,
                 reg1235,
                 reg1230,
                 reg1229,
                 reg1226,
                 reg1223,
                 reg1222,
                 reg1219,
                 reg1218,
                 reg1217,
                 reg1214,
                 reg1213,
                 reg1210,
                 reg1209,
                 reg1207,
                 reg1205,
                 reg1204,
                 reg1199,
                 reg1200,
                 reg1286,
                 reg1285,
                 reg1281,
                 reg1279,
                 reg1277,
                 reg1275,
                 reg1274,
                 reg1273,
                 reg1272,
                 reg1271,
                 reg1270,
                 reg1269,
                 reg1268,
                 reg1267,
                 reg1264,
                 reg1262,
                 reg1261,
                 reg1260,
                 reg1259,
                 reg1256,
                 forvar1255,
                 reg1252,
                 reg1247,
                 reg1244,
                 reg1242,
                 reg1241,
                 reg1240,
                 reg1239,
                 forvar1237,
                 reg1236,
                 reg1234,
                 reg1233,
                 forvar1232,
                 reg1231,
                 reg1228,
                 forvar1227,
                 reg1225,
                 reg1224,
                 forvar1221,
                 reg1220,
                 forvar1216,
                 reg1215,
                 reg1208,
                 reg1206,
                 reg1203,
                 reg1202,
                 reg1201,
                 forvar1199,
                 reg1198,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned(wire1195[(5'h11):(3'h4)]))
        begin
          reg1198 = $signed(wire1194);
          for (forvar1199 = (1'h0); (forvar1199 < (1'h0)); forvar1199 = (forvar1199 + (1'h1)))
            begin
              reg1200 <= (wire1195 & ({wire1193,
                      ((wire1194 ? wire1193 : wire1193) ?
                          $unsigned(wire1193) : $unsigned(wire1194))} ?
                  reg1198[(3'h5):(1'h1)] : ($unsigned(wire1193) * $signed(wire1195))));
              reg1201 = $signed((~&$signed((wire1196[(4'h9):(3'h7)] ?
                  (8'ha4) : (forvar1199 ? reg1200 : wire1194)))));
              reg1202 = (wire1194 ? $unsigned(wire1195) : wire1196);
            end
        end
      else
        begin
          reg1198 = ((7'h48) ?
              ({reg1201[(4'h8):(3'h6)], ((|reg1201) | ((7'h44) ~^ reg1200))} ?
                  reg1202[(4'hc):(4'ha)] : wire1195[(2'h3):(2'h3)]) : (+(^~((8'hb3) ?
                  $signed(reg1201) : (wire1195 ? wire1195 : wire1193)))));
          if ($signed(wire1194[(1'h0):(1'h0)]))
            begin
              reg1199 <= $signed($signed(wire1193));
            end
          else
            begin
              reg1201 = (wire1196[(4'h8):(2'h3)] && wire1194);
              reg1202 = wire1197[(5'h12):(2'h3)];
              reg1203 = ((wire1195[(4'hf):(3'h4)] - ($signed(reg1200) ?
                      (-(forvar1199 <= reg1201)) : $signed((wire1197 + wire1194)))) ?
                  $signed(reg1198) : ({($signed(wire1195) <= (wire1193 ?
                              reg1201 : reg1202)),
                          ((^~reg1198) ?
                              (wire1196 ?
                                  wire1195 : wire1194) : (wire1193 == wire1195))} ?
                      reg1200[(1'h1):(1'h1)] : (|(wire1194[(5'h16):(5'h13)] ?
                          reg1198[(4'h8):(2'h3)] : wire1197))));
            end
          if ((wire1196[(3'h7):(2'h2)] | ($unsigned($signed({reg1199,
              (7'h49)})) * (forvar1199[(3'h6):(1'h1)] & {$signed(reg1199)}))))
            begin
              reg1204 <= $signed(({{(reg1202 ? (8'ha7) : forvar1199),
                      (wire1195 <= reg1202)},
                  $signed((wire1193 ^ wire1193))} | $unsigned(reg1200)));
              reg1205 <= (wire1193[(3'h6):(1'h0)] ~^ reg1200);
              reg1206 = ((wire1193[(3'h6):(1'h0)] + $unsigned(($unsigned(reg1200) ?
                      $signed(reg1198) : (+reg1198)))) ?
                  {((&$signed(reg1202)) ?
                          {$signed((8'hb0))} : $signed((reg1202 ?
                              (8'h9d) : reg1203))),
                      {$signed(((8'ha1) ^~ reg1200))}} : (~&$signed($unsigned($signed(wire1194)))));
            end
          else
            begin
              reg1204 <= $signed((^~((reg1204 << wire1197[(3'h6):(2'h3)]) ?
                  reg1202[(3'h6):(3'h4)] : ((reg1201 ? forvar1199 : (8'h9c)) ?
                      forvar1199[(3'h5):(1'h1)] : (reg1200 == reg1204)))));
            end
          if ((reg1203 >>> reg1198[(4'h9):(3'h5)]))
            begin
              reg1207 <= $signed({((~(reg1204 ? reg1202 : wire1196)) ?
                      $unsigned((wire1193 ? reg1206 : reg1201)) : (7'h43)),
                  (~|(reg1204[(2'h3):(1'h1)] | {wire1197, reg1205}))});
            end
          else
            begin
              reg1208 = $unsigned(reg1198[(3'h6):(3'h4)]);
            end
          reg1209 <= (~&((+reg1206[(3'h5):(1'h1)]) ?
              reg1204[(4'hf):(1'h1)] : ((|((8'hbd) >> wire1197)) ?
                  $signed((reg1199 ? (8'ha6) : reg1199)) : ((reg1206 ?
                          forvar1199 : wire1195) ?
                      reg1207[(4'hc):(4'hc)] : reg1206))));
        end
      reg1210 <= ((+(($signed((8'hb0)) ^ reg1206[(3'h5):(3'h4)]) ?
              ($signed(wire1193) ?
                  {(8'hb9), wire1194} : $unsigned(reg1209)) : (7'h47))) ?
          reg1203[(1'h0):(1'h0)] : $unsigned((({wire1193} ?
                  (reg1205 ? (8'hae) : reg1205) : reg1203[(4'hf):(4'hb)]) ?
              $unsigned(forvar1199) : reg1207)));
    end
  assign wire1211 = (~&reg1205);
  assign wire1212 = $signed($signed($unsigned(wire1195[(4'he):(2'h3)])));
  always
    @(posedge clk) begin
      reg1213 <= (^wire1194);
      reg1214 <= reg1213;
      reg1215 = reg1204;
      for (forvar1216 = (1'h0); (forvar1216 < (2'h2)); forvar1216 = (forvar1216 + (1'h1)))
        begin
          reg1217 <= (~&((({(8'hb7)} > {reg1215}) ^~ $unsigned(reg1215[(1'h1):(1'h0)])) ?
              wire1197 : reg1215[(3'h4):(3'h4)]));
          reg1218 <= ({{($signed(wire1194) ? (reg1204 >> wire1212) : wire1211),
                  reg1207[(5'h10):(4'hf)]},
              $signed(($signed(reg1214) == (reg1200 + reg1205)))} >> ({$signed((~&wire1197)),
              ((+wire1195) ? (wire1197 ^ wire1197) : reg1200)} < (((reg1207 ?
                      wire1212 : (7'h4a)) ?
                  $unsigned((8'hb6)) : wire1193[(4'h9):(2'h3)]) ?
              $unsigned($signed(forvar1216)) : reg1207[(4'hc):(4'h9)])));
          reg1219 <= $unsigned(reg1209);
          reg1220 = (reg1214[(1'h1):(1'h0)] ? (8'ha9) : wire1194);
          for (forvar1221 = (1'h0); (forvar1221 < (1'h1)); forvar1221 = (forvar1221 + (1'h1)))
            begin
              reg1222 <= ((8'haf) ^~ ((!reg1213[(3'h7):(3'h7)]) ?
                  $signed((((8'haf) ?
                      reg1205 : (8'hb5)) >>> reg1217[(2'h2):(1'h1)])) : reg1218[(3'h4):(2'h2)]));
              reg1223 <= (~(!(|(8'hbe))));
              reg1224 = reg1218[(4'hc):(1'h1)];
              reg1225 = reg1214[(4'h8):(1'h0)];
              reg1226 <= (^~((~|reg1199[(1'h0):(1'h0)]) ?
                  $signed($signed(reg1219[(3'h6):(2'h3)])) : ((+$unsigned(wire1195)) * {$unsigned(wire1195),
                      $unsigned(reg1214)})));
            end
        end
      if ($unsigned((&(((|reg1224) > (reg1219 ?
          wire1193 : reg1204)) && $unsigned((reg1209 ? reg1220 : wire1193))))))
        begin
          for (forvar1227 = (1'h0); (forvar1227 < (3'h4)); forvar1227 = (forvar1227 + (1'h1)))
            begin
              reg1228 = forvar1216[(4'hb):(4'ha)];
            end
        end
      else
        begin
          for (forvar1227 = (1'h0); (forvar1227 < (1'h0)); forvar1227 = (forvar1227 + (1'h1)))
            begin
              reg1228 = (8'ha2);
              reg1229 <= (~(^wire1212));
              reg1230 <= wire1197;
            end
        end
    end
  always
    @(posedge clk) begin
      reg1231 = ($signed(reg1219) ^~ {wire1194,
          ($signed($signed(wire1194)) ^ (wire1211 ^~ wire1212))});
      for (forvar1232 = (1'h0); (forvar1232 < (1'h0)); forvar1232 = (forvar1232 + (1'h1)))
        begin
          if (({wire1211[(2'h2):(1'h0)]} ?
              $signed(reg1210[(1'h0):(1'h0)]) : (reg1204[(2'h3):(2'h3)] == reg1231)))
            begin
              reg1233 = (&$signed($signed(reg1200)));
            end
          else
            begin
              reg1233 = (!reg1223);
              reg1234 = (~|(wire1194[(4'hd):(4'hc)] << $signed($signed(((8'hbb) ?
                  reg1205 : (8'hb3))))));
            end
          if ($signed(($signed((~&(|wire1194))) > $signed(($signed(reg1226) & (reg1199 ?
              (8'hac) : (7'h45)))))))
            begin
              reg1235 <= (((+reg1218[(3'h7):(3'h6)]) ?
                      ($unsigned((wire1212 ^~ wire1196)) ?
                          reg1219 : $signed((^(8'hb2)))) : reg1204) ?
                  (!$signed($signed((7'h42)))) : $unsigned((|$unsigned($signed(reg1234)))));
            end
          else
            begin
              reg1235 <= ($signed((($unsigned(forvar1232) >> reg1207[(4'hf):(2'h3)]) >= (^~((7'h43) && reg1235)))) <= (-$unsigned(((reg1199 <= wire1212) ~^ (wire1196 <= reg1231)))));
            end
          reg1236 = reg1230[(4'hc):(4'h8)];
          for (forvar1237 = (1'h0); (forvar1237 < (1'h1)); forvar1237 = (forvar1237 + (1'h1)))
            begin
              reg1238 <= ($signed(reg1226[(2'h3):(1'h1)]) != (($unsigned((reg1234 ^~ reg1222)) <<< reg1236) != $signed($signed(wire1196[(4'hb):(4'h8)]))));
              reg1239 = (~reg1214);
              reg1240 = {$signed(({((8'hac) << wire1212),
                      forvar1237} ^ ($signed(reg1217) ?
                      reg1226[(3'h6):(1'h1)] : reg1234[(4'hd):(4'h9)]))),
                  ($unsigned((7'h42)) ?
                      $signed((!reg1226)) : {(^~(!(8'ha4)))})};
            end
          if ((reg1217 * wire1212[(3'h5):(3'h4)]))
            begin
              reg1241 = reg1240[(3'h6):(1'h1)];
            end
          else
            begin
              reg1241 = reg1205;
            end
        end
      reg1242 = reg1213;
      if (wire1194)
        begin
          if ((~$signed(reg1236[(3'h6):(2'h2)])))
            begin
              reg1243 <= reg1236[(3'h7):(3'h7)];
              reg1244 = wire1194[(4'h9):(4'h9)];
              reg1245 <= reg1241;
              reg1246 <= (^$unsigned((!$signed($unsigned(wire1194)))));
            end
          else
            begin
              reg1244 = ((~&wire1193) * ((reg1209 ?
                      $unsigned({wire1211, reg1239}) : (!((8'hb2) ?
                          reg1235 : reg1246))) ?
                  (8'hb8) : $signed(($signed(wire1212) ?
                      (forvar1237 || wire1194) : $signed(wire1195)))));
              reg1245 <= reg1205[(4'hc):(1'h1)];
              reg1246 <= reg1226[(2'h2):(1'h1)];
              reg1247 = (!$unsigned(reg1209));
              reg1248 <= (8'ha3);
            end
          if ($unsigned($signed((8'hab))))
            begin
              reg1249 <= (!(($unsigned(reg1248) ?
                  (~^reg1222) : $unsigned($unsigned(reg1248))) >>> reg1245[(2'h2):(1'h0)]));
              reg1250 <= ((reg1230[(3'h5):(1'h0)] ^ ((&$signed(reg1205)) ?
                  wire1197 : (~&((7'h48) ?
                      wire1194 : reg1204)))) <<< (($unsigned((~&(8'ha2))) <<< (!$unsigned(reg1239))) * $signed(reg1222)));
              reg1251 <= reg1205[(4'hb):(1'h0)];
              reg1252 = $unsigned(($signed((8'hb0)) & (~^($unsigned((7'h42)) && $signed(reg1217)))));
              reg1253 <= $signed(forvar1232);
            end
          else
            begin
              reg1249 <= reg1209;
            end
          reg1254 <= reg1248[(4'h9):(4'h8)];
          for (forvar1255 = (1'h0); (forvar1255 < (3'h4)); forvar1255 = (forvar1255 + (1'h1)))
            begin
              reg1256 = reg1204[(5'h11):(4'h8)];
              reg1257 <= reg1204[(1'h1):(1'h1)];
              reg1258 <= (8'hb3);
            end
          reg1259 = (+forvar1232[(3'h7):(3'h7)]);
        end
      else
        begin
          reg1244 = reg1251[(3'h4):(1'h1)];
        end
      if (reg1253[(4'hd):(4'ha)])
        begin
          reg1260 = (~{(~(~|$signed(reg1241))), (~^{reg1253[(5'h13):(4'h8)]})});
          if ({forvar1255, $signed(reg1259)})
            begin
              reg1261 = ({$signed(reg1252[(2'h2):(1'h1)])} ?
                  (^~(+($signed((8'hab)) ?
                      (reg1254 ^~ reg1205) : $unsigned(reg1209)))) : $signed(reg1236[(2'h3):(1'h1)]));
              reg1262 = (((reg1209 <= $signed($signed(reg1219))) == reg1253) == wire1197);
              reg1263 <= $unsigned((!$signed((^(^~reg1258)))));
            end
          else
            begin
              reg1263 <= (reg1239[(3'h4):(2'h2)] && $signed($signed({reg1246[(4'he):(3'h6)],
                  ((8'ha4) ? reg1263 : reg1240)})));
            end
          if (wire1195)
            begin
              reg1264 = ({reg1235,
                  ($signed($unsigned((8'hb0))) ?
                      $unsigned((reg1229 != reg1200)) : $unsigned(((7'h46) ^ wire1195)))} ^ {($signed((reg1247 ?
                      reg1229 : wire1193)) & $signed($unsigned(reg1258)))});
              reg1265 <= reg1264[(3'h4):(1'h1)];
              reg1266 <= reg1246;
              reg1267 = reg1250;
            end
          else
            begin
              reg1264 = reg1249[(4'hb):(3'h5)];
              reg1267 = {$signed((|$unsigned(reg1238)))};
              reg1268 = reg1209;
              reg1269 = reg1222;
              reg1270 = (+{$unsigned((~^(8'hac)))});
            end
          if (((!reg1213[(2'h3):(2'h2)]) ?
              (^{$unsigned((reg1226 | (8'haa)))}) : $unsigned((({wire1193,
                      (8'hb9)} ^ (reg1240 ? reg1267 : reg1265)) ?
                  forvar1232 : (reg1213[(2'h2):(1'h0)] ?
                      {reg1266, (8'hb2)} : reg1243[(3'h4):(2'h3)])))))
            begin
              reg1271 = (reg1236[(4'ha):(4'h9)] >= $signed($unsigned({$unsigned(reg1246),
                  ((8'hb7) ^~ reg1199)})));
              reg1272 = forvar1237;
              reg1273 = (&$signed((reg1235[(1'h1):(1'h0)] ~^ ((-reg1207) ?
                  {(8'hb9)} : (!reg1258)))));
              reg1274 = $signed(reg1235[(4'hc):(3'h7)]);
              reg1275 = ((^(~(reg1242 < reg1241))) != forvar1232);
            end
          else
            begin
              reg1276 <= $unsigned(reg1214[(4'h9):(3'h5)]);
              reg1277 = {((($signed((8'h9d)) < reg1266[(2'h3):(2'h3)]) + (!$signed((8'h9c)))) ?
                      reg1209[(4'h9):(4'h9)] : reg1259)};
              reg1278 <= reg1251[(1'h1):(1'h0)];
              reg1279 = reg1252;
            end
          if ({reg1252, (~|(~^(8'hbe)))})
            begin
              reg1280 <= ($signed(((!(^reg1249)) ~^ forvar1232[(2'h2):(1'h1)])) ?
                  {(+((8'ha1) * reg1278)),
                      ($signed($signed(reg1262)) != {(reg1205 ?
                              (8'ha8) : reg1270),
                          reg1199[(4'h8):(3'h6)]})} : $unsigned($unsigned({$unsigned(reg1259),
                      $unsigned(reg1207)})));
              reg1281 = reg1231;
              reg1282 <= (~&(($signed((&reg1281)) * $signed((^~reg1263))) == reg1214[(4'hc):(4'h8)]));
              reg1283 <= reg1249[(3'h6):(2'h2)];
              reg1284 <= $unsigned(({(reg1230[(4'hb):(1'h0)] ?
                          (reg1268 <<< reg1272) : $signed(reg1252))} ?
                  ($unsigned((reg1233 ? reg1233 : (8'h9f))) ?
                      (-$signed(reg1233)) : $signed($signed(reg1222))) : $signed($signed((~^reg1229)))));
            end
          else
            begin
              reg1280 <= reg1284[(5'h11):(2'h2)];
              reg1281 = $unsigned(($unsigned($unsigned(reg1265)) * $unsigned((reg1271[(4'hd):(3'h5)] * $signed((8'had))))));
              reg1282 <= {$signed(reg1248[(1'h1):(1'h1)]),
                  (|$unsigned(reg1234))};
              reg1285 = $signed((^(reg1241[(1'h1):(1'h0)] & ((8'ha7) ~^ reg1239[(3'h4):(2'h2)]))));
              reg1286 = $unsigned(reg1217[(4'h8):(1'h1)]);
            end
        end
      else
        begin
          if ((~^($unsigned((+(reg1249 ? wire1211 : reg1257))) >>> {({reg1283,
                  reg1200} & forvar1232)})))
            begin
              reg1260 = ({reg1272[(3'h5):(2'h2)]} + $unsigned((~|($unsigned(reg1209) >>> $signed(wire1195)))));
              reg1263 <= $unsigned(($signed({$signed(reg1200),
                  ((8'hb4) ? reg1248 : (8'ha6))}) >>> {((reg1229 == reg1279) ?
                      (8'hbe) : $unsigned(reg1274)),
                  ({reg1243} + {reg1279, reg1284})}));
              reg1264 = (^(7'h48));
              reg1265 <= reg1243[(2'h2):(2'h2)];
              reg1266 <= {reg1261, (8'ha6)};
            end
          else
            begin
              reg1260 = (^(($signed(reg1219) ?
                      ((reg1270 ?
                          reg1223 : (8'hb9)) ~^ (~^(8'hb2))) : ((+reg1199) ?
                          $unsigned((8'hb3)) : (reg1223 < reg1263))) ?
                  (^{reg1271}) : {((wire1194 ? reg1205 : (8'hb6)) ?
                          (reg1213 | reg1279) : (reg1231 ?
                              wire1195 : wire1193)),
                      (8'h9f)}));
              reg1261 = {((-reg1246) ?
                      $unsigned(reg1236) : (+reg1286[(4'h8):(2'h3)])),
                  reg1241[(5'h15):(3'h5)]};
              reg1263 <= $signed({$signed($signed((reg1276 ?
                      reg1210 : reg1282)))});
              reg1264 = reg1200[(1'h1):(1'h0)];
            end
          reg1276 <= wire1197;
          if (reg1207)
            begin
              reg1277 = $unsigned($unsigned(({wire1196[(1'h1):(1'h1)]} ?
                  $unsigned((reg1262 ?
                      (7'h49) : (8'ha0))) : (reg1240[(3'h7):(3'h5)] & $unsigned(reg1261)))));
              reg1278 <= reg1241;
              reg1280 <= (&reg1247);
            end
          else
            begin
              reg1277 = reg1233[(2'h2):(1'h0)];
              reg1279 = reg1259[(2'h2):(1'h0)];
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module1025  (y, clk, wire1030, wire1029, wire1028, wire1027, wire1026);
  output wire [(32'h7c4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire1030;
  input wire signed [(5'h15):(1'h0)] wire1029;
  input wire [(3'h6):(1'h0)] wire1028;
  input wire [(4'hd):(1'h0)] wire1027;
  input wire [(3'h5):(1'h0)] wire1026;
  wire signed [(3'h6):(1'h0)] wire1138;
  wire signed [(4'he):(1'h0)] wire1126;
  wire signed [(5'h11):(1'h0)] wire1125;
  wire signed [(2'h2):(1'h0)] wire1124;
  wire [(4'hb):(1'h0)] wire1123;
  wire signed [(5'h10):(1'h0)] wire1122;
  wire [(4'hd):(1'h0)] wire1121;
  wire [(5'h17):(1'h0)] wire1120;
  wire signed [(5'h14):(1'h0)] wire1054;
  wire [(4'h9):(1'h0)] wire1053;
  reg signed [(5'h17):(1'h0)] reg1166 = (1'h0);
  reg [(5'h15):(1'h0)] reg1164 = (1'h0);
  reg [(3'h4):(1'h0)] reg1163 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1161 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1153 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1152 = (1'h0);
  reg [(4'hc):(1'h0)] reg1150 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1146 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1144 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1141 = (1'h0);
  reg [(5'h14):(1'h0)] reg1137 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1133 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1131 = (1'h0);
  reg [(5'h16):(1'h0)] reg1127 = (1'h0);
  reg [(2'h2):(1'h0)] reg1119 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1118 = (1'h0);
  reg [(5'h13):(1'h0)] reg1114 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1116 = (1'h0);
  reg [(5'h17):(1'h0)] reg1105 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1103 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1099 = (1'h0);
  reg [(2'h2):(1'h0)] reg1097 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1092 = (1'h0);
  reg [(5'h17):(1'h0)] reg1096 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1094 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1090 = (1'h0);
  reg [(4'h8):(1'h0)] reg1087 = (1'h0);
  reg [(2'h3):(1'h0)] reg1086 = (1'h0);
  reg [(4'hc):(1'h0)] reg1083 = (1'h0);
  reg [(4'h9):(1'h0)] reg1076 = (1'h0);
  reg [(3'h6):(1'h0)] reg1074 = (1'h0);
  reg [(5'h11):(1'h0)] reg1073 = (1'h0);
  reg [(5'h10):(1'h0)] reg1067 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1064 = (1'h0);
  reg [(4'h8):(1'h0)] reg1063 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1062 = (1'h0);
  reg [(4'hd):(1'h0)] reg1057 = (1'h0);
  reg [(4'hd):(1'h0)] reg1055 = (1'h0);
  reg [(5'h10):(1'h0)] reg1052 = (1'h0);
  reg [(5'h16):(1'h0)] reg1051 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1049 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1047 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1046 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1045 = (1'h0);
  reg [(3'h5):(1'h0)] reg1041 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1039 = (1'h0);
  reg [(4'ha):(1'h0)] reg1038 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1036 = (1'h0);
  reg [(5'h11):(1'h0)] reg1035 = (1'h0);
  reg [(5'h17):(1'h0)] reg1034 = (1'h0);
  reg [(5'h10):(1'h0)] reg1032 = (1'h0);
  reg [(2'h3):(1'h0)] reg1165 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1162 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1160 = (1'h0);
  reg [(5'h17):(1'h0)] reg1159 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1158 = (1'h0);
  reg [(5'h11):(1'h0)] reg1157 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1156 = (1'h0);
  reg [(4'h9):(1'h0)] reg1155 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1154 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1151 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1149 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1148 = (1'h0);
  reg [(5'h11):(1'h0)] reg1147 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1145 = (1'h0);
  reg [(3'h5):(1'h0)] forvar1143 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1142 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar1140 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1139 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1136 = (1'h0);
  reg [(4'he):(1'h0)] reg1135 = (1'h0);
  reg [(5'h15):(1'h0)] reg1134 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1133 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1127 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1132 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1130 = (1'h0);
  reg [(4'hb):(1'h0)] reg1129 = (1'h0);
  reg [(5'h10):(1'h0)] reg1128 = (1'h0);
  reg [(4'h9):(1'h0)] reg1109 = (1'h0);
  reg [(5'h13):(1'h0)] reg1117 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1115 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1114 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1113 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1112 = (1'h0);
  reg [(3'h5):(1'h0)] reg1111 = (1'h0);
  reg [(4'hc):(1'h0)] reg1110 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar1109 = (1'h0);
  reg [(3'h4):(1'h0)] reg1108 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1107 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1106 = (1'h0);
  reg [(3'h5):(1'h0)] reg1104 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1102 = (1'h0);
  reg [(2'h2):(1'h0)] reg1101 = (1'h0);
  reg [(3'h5):(1'h0)] reg1100 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1098 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1087 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1095 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1093 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1092 = (1'h0);
  reg [(4'h8):(1'h0)] reg1091 = (1'h0);
  reg [(4'h9):(1'h0)] reg1089 = (1'h0);
  reg [(2'h2):(1'h0)] reg1088 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1080 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1085 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1084 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1082 = (1'h0);
  reg [(5'h17):(1'h0)] reg1081 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1080 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1079 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1078 = (1'h0);
  reg [(2'h3):(1'h0)] reg1077 = (1'h0);
  reg [(5'h16):(1'h0)] reg1075 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1073 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1071 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1067 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1072 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar1071 = (1'h0);
  reg [(3'h4):(1'h0)] reg1070 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1069 = (1'h0);
  reg [(5'h11):(1'h0)] reg1068 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1066 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1065 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1061 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1060 = (1'h0);
  reg [(4'he):(1'h0)] reg1059 = (1'h0);
  reg [(5'h18):(1'h0)] reg1058 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1056 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar1055 = (1'h0);
  reg [(5'h17):(1'h0)] reg1050 = (1'h0);
  reg [(4'ha):(1'h0)] reg1048 = (1'h0);
  reg [(5'h15):(1'h0)] reg1044 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1043 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1042 = (1'h0);
  reg [(5'h11):(1'h0)] reg1040 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1033 = (1'h0);
  reg [(5'h15):(1'h0)] reg1037 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1033 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1031 = (1'h0);
  assign y = {wire1138,
                 wire1126,
                 wire1125,
                 wire1124,
                 wire1123,
                 wire1122,
                 wire1121,
                 wire1120,
                 wire1054,
                 wire1053,
                 reg1166,
                 reg1164,
                 reg1163,
                 reg1161,
                 reg1153,
                 reg1152,
                 reg1150,
                 reg1146,
                 reg1144,
                 reg1141,
                 reg1137,
                 reg1133,
                 reg1131,
                 reg1127,
                 reg1119,
                 reg1118,
                 reg1114,
                 reg1116,
                 reg1105,
                 reg1103,
                 reg1099,
                 reg1097,
                 reg1092,
                 reg1096,
                 reg1094,
                 reg1090,
                 reg1087,
                 reg1086,
                 reg1083,
                 reg1076,
                 reg1074,
                 reg1073,
                 reg1067,
                 reg1064,
                 reg1063,
                 reg1062,
                 reg1057,
                 reg1055,
                 reg1052,
                 reg1051,
                 reg1049,
                 reg1047,
                 reg1046,
                 reg1045,
                 reg1041,
                 reg1039,
                 reg1038,
                 reg1036,
                 reg1035,
                 reg1034,
                 reg1032,
                 reg1165,
                 reg1162,
                 forvar1160,
                 reg1159,
                 reg1158,
                 reg1157,
                 reg1156,
                 reg1155,
                 forvar1154,
                 reg1151,
                 reg1149,
                 forvar1148,
                 reg1147,
                 reg1145,
                 forvar1143,
                 reg1142,
                 forvar1140,
                 forvar1139,
                 reg1136,
                 reg1135,
                 reg1134,
                 forvar1133,
                 forvar1127,
                 reg1132,
                 reg1130,
                 reg1129,
                 reg1128,
                 reg1109,
                 reg1117,
                 reg1115,
                 forvar1114,
                 reg1113,
                 reg1112,
                 reg1111,
                 reg1110,
                 forvar1109,
                 reg1108,
                 reg1107,
                 forvar1106,
                 reg1104,
                 reg1102,
                 reg1101,
                 reg1100,
                 forvar1098,
                 forvar1087,
                 reg1095,
                 reg1093,
                 forvar1092,
                 reg1091,
                 reg1089,
                 reg1088,
                 forvar1080,
                 reg1085,
                 reg1084,
                 reg1082,
                 reg1081,
                 reg1080,
                 reg1079,
                 reg1078,
                 reg1077,
                 reg1075,
                 forvar1073,
                 reg1071,
                 forvar1067,
                 reg1072,
                 forvar1071,
                 reg1070,
                 reg1069,
                 reg1068,
                 reg1066,
                 reg1065,
                 forvar1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 reg1056,
                 forvar1055,
                 reg1050,
                 reg1048,
                 reg1044,
                 reg1043,
                 forvar1042,
                 reg1040,
                 forvar1033,
                 reg1037,
                 reg1033,
                 reg1031,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg1031 = wire1028[(3'h5):(2'h2)];
      reg1032 <= wire1027[(2'h2):(1'h0)];
      if (((wire1028 ?
              ((wire1029[(4'h9):(3'h5)] & $signed(wire1029)) ?
                  (reg1032[(3'h5):(3'h5)] ?
                      $unsigned(wire1030) : $unsigned(wire1028)) : (~$signed((8'hbf)))) : (^~wire1028)) ?
          $unsigned(wire1029[(3'h4):(3'h4)]) : (+wire1028[(3'h4):(1'h1)])))
        begin
          if ((8'hbe))
            begin
              reg1033 = $unsigned(($unsigned(({wire1028, wire1026} ?
                  wire1030[(1'h0):(1'h0)] : $signed(wire1028))) == $unsigned(({reg1032} <<< (reg1031 ?
                  reg1032 : reg1032)))));
              reg1034 <= ($unsigned(($signed((^wire1026)) ?
                      ({reg1031} ?
                          (reg1031 ?
                              reg1031 : wire1030) : $unsigned((7'h40))) : {(wire1029 ?
                              reg1031 : wire1030)})) ?
                  wire1028[(1'h0):(1'h0)] : $unsigned($signed(((wire1028 ?
                          reg1033 : wire1030) ?
                      (+wire1029) : (reg1033 ? wire1026 : reg1033)))));
              reg1035 <= $unsigned({(8'h9d)});
            end
          else
            begin
              reg1034 <= (-{$unsigned((reg1033[(4'h9):(3'h4)] && (wire1030 ?
                      reg1032 : (8'hab)))),
                  wire1026});
              reg1035 <= reg1035[(5'h11):(4'hd)];
              reg1036 <= $unsigned((|($signed($unsigned(reg1032)) == $signed((~reg1032)))));
              reg1037 = $signed(({($signed(reg1036) << (reg1031 ?
                      wire1028 : wire1030)),
                  $signed($signed(wire1026))} + reg1036[(2'h2):(2'h2)]));
              reg1038 <= (reg1031[(3'h7):(2'h2)] ^~ reg1031);
            end
          reg1039 <= wire1026;
        end
      else
        begin
          for (forvar1033 = (1'h0); (forvar1033 < (1'h1)); forvar1033 = (forvar1033 + (1'h1)))
            begin
              reg1037 = $unsigned($signed($unsigned((-(8'hac)))));
            end
          if (wire1030[(1'h1):(1'h0)])
            begin
              reg1040 = wire1029[(4'h9):(2'h2)];
            end
          else
            begin
              reg1038 <= (~{reg1034});
              reg1039 <= (~&$unsigned((reg1038[(4'h8):(1'h0)] ?
                  {(~reg1038), $signed(reg1040)} : (+(~&reg1040)))));
              reg1041 <= $unsigned(($unsigned(((~^(8'h9d)) ?
                      (^~wire1030) : (wire1026 >= reg1035))) ?
                  {$signed((forvar1033 ?
                          reg1034 : wire1027))} : (reg1037[(4'h8):(4'h8)] ?
                      wire1029[(4'hf):(4'hc)] : ((forvar1033 ?
                              reg1037 : reg1032) ?
                          $signed(wire1028) : $unsigned(reg1036)))));
            end
          for (forvar1042 = (1'h0); (forvar1042 < (1'h0)); forvar1042 = (forvar1042 + (1'h1)))
            begin
              reg1043 = wire1028[(3'h6):(3'h5)];
              reg1044 = $unsigned($signed($unsigned(((reg1039 ?
                  forvar1033 : reg1040) <<< (reg1039 ? reg1033 : reg1037)))));
              reg1045 <= (~(|($unsigned((reg1031 + reg1032)) >> ($unsigned(reg1033) ?
                  reg1037[(4'hf):(2'h3)] : reg1041))));
              reg1046 <= reg1041[(3'h4):(2'h2)];
              reg1047 <= $unsigned(({{$signed(reg1044)}} ?
                  wire1030 : $unsigned($unsigned(reg1037))));
            end
          if (reg1035[(1'h1):(1'h1)])
            begin
              reg1048 = {reg1043[(4'hd):(3'h6)]};
              reg1049 <= ((&((7'h43) ?
                  (&$unsigned(reg1037)) : $unsigned(reg1041))) < (~$unsigned($signed((reg1041 << wire1028)))));
              reg1050 = ($unsigned((~&{(reg1044 ^~ reg1047),
                  (reg1031 >= reg1031)})) <<< $unsigned({reg1043[(4'he):(4'he)]}));
            end
          else
            begin
              reg1049 <= reg1036[(2'h2):(1'h1)];
              reg1050 = $unsigned({((+(reg1037 && reg1047)) ^~ reg1039),
                  $signed(wire1030[(1'h0):(1'h0)])});
              reg1051 <= $signed(reg1039);
            end
        end
      reg1052 <= $signed((7'h41));
    end
  assign wire1053 = (&(($signed((^reg1046)) ?
                        reg1049 : reg1047[(4'he):(3'h4)]) + (reg1038[(3'h5):(1'h1)] ?
                        reg1038 : (-reg1049[(5'h14):(5'h14)]))));
  assign wire1054 = $unsigned(($signed(reg1045[(4'hf):(4'hb)]) + ((-(wire1053 <= (7'h43))) ?
                        $signed((reg1038 + reg1045)) : (|wire1026[(1'h1):(1'h1)]))));
  always
    @(posedge clk) begin
      if (({(8'hbe)} ?
          (~^({reg1051[(3'h5):(2'h3)]} ?
              (wire1026 <= reg1052) : reg1051[(2'h2):(1'h1)])) : ((~^({reg1047} >> (reg1051 ~^ wire1054))) | (($unsigned((7'h41)) <<< (wire1030 ?
              reg1051 : reg1032)) == ((~^wire1029) ?
              $signed(wire1028) : $unsigned(reg1049))))))
        begin
          for (forvar1055 = (1'h0); (forvar1055 < (3'h4)); forvar1055 = (forvar1055 + (1'h1)))
            begin
              reg1056 = reg1049[(4'hc):(3'h6)];
            end
        end
      else
        begin
          if (reg1034)
            begin
              reg1055 <= (~|((reg1034[(4'he):(3'h6)] ?
                      ($signed(reg1051) ?
                          (reg1047 * reg1038) : reg1051) : $signed((8'ha5))) ?
                  (wire1029[(5'h15):(4'hc)] ?
                      ($unsigned(wire1029) ?
                          $signed(reg1047) : wire1028[(3'h5):(3'h4)]) : $unsigned({reg1052,
                          wire1030})) : {(reg1051[(5'h15):(3'h4)] && (-wire1026))}));
              reg1056 = (wire1054 * $unsigned($unsigned(wire1054[(2'h2):(1'h0)])));
              reg1057 <= wire1027;
              reg1058 = (wire1053[(1'h0):(1'h0)] >= $signed(($signed($unsigned(wire1028)) - {reg1045,
                  (reg1055 ? wire1028 : reg1057)})));
            end
          else
            begin
              reg1056 = $signed({$unsigned((reg1056 + (wire1029 || reg1035))),
                  ({$unsigned(forvar1055), reg1035} ?
                      $signed($signed(reg1034)) : ((~^reg1038) ^ (~^(8'ha4))))});
              reg1058 = (~&reg1047[(3'h5):(1'h1)]);
            end
          reg1059 = (~^((&wire1028[(3'h4):(2'h3)]) <<< (wire1026[(2'h2):(1'h0)] ?
              (7'h42) : wire1054)));
          reg1060 = reg1058[(3'h4):(3'h4)];
          for (forvar1061 = (1'h0); (forvar1061 < (1'h0)); forvar1061 = (forvar1061 + (1'h1)))
            begin
              reg1062 <= (!(!($signed($signed(reg1045)) >= ((reg1059 ?
                      reg1034 : forvar1055) ?
                  (wire1053 != reg1036) : forvar1061))));
              reg1063 <= (wire1027[(4'hc):(3'h5)] * wire1029[(3'h6):(1'h1)]);
            end
          reg1064 <= wire1029;
        end
      reg1065 = reg1046;
      reg1066 = ($signed(reg1036) ?
          $unsigned(($unsigned((reg1062 <<< reg1062)) >= $signed((8'ha9)))) : ((~(reg1058 ?
              $unsigned(wire1028) : reg1060)) | {$signed((~&wire1030)),
              $unsigned($signed(reg1055))}));
      if (wire1054[(5'h12):(3'h7)])
        begin
          reg1067 <= (($unsigned($signed((^~wire1029))) - $unsigned((~|(reg1045 ?
              wire1030 : forvar1061)))) * {reg1055,
              $signed((reg1066[(2'h3):(2'h2)] ?
                  (^reg1063) : $signed(reg1052)))});
          reg1068 = $unsigned((-reg1032));
          reg1069 = {{reg1065, wire1026}, forvar1055[(5'h12):(1'h0)]};
          reg1070 = (reg1068[(3'h5):(1'h0)] ?
              ((wire1054 <= (reg1032 + (reg1057 ~^ (8'ha3)))) <<< ($unsigned((wire1030 ?
                  (8'ha1) : reg1062)) >> reg1055)) : $unsigned($signed((~^(reg1045 || reg1036)))));
          for (forvar1071 = (1'h0); (forvar1071 < (2'h2)); forvar1071 = (forvar1071 + (1'h1)))
            begin
              reg1072 = $signed((&$unsigned((^~(reg1046 || reg1045)))));
              reg1073 <= wire1026;
              reg1074 <= {reg1069,
                  ((!reg1070[(2'h2):(1'h1)]) ?
                      $unsigned((reg1055 ?
                          (forvar1055 ? reg1069 : reg1052) : (reg1070 ?
                              reg1066 : reg1051))) : (-$signed((&reg1066))))};
            end
        end
      else
        begin
          for (forvar1067 = (1'h0); (forvar1067 < (1'h1)); forvar1067 = (forvar1067 + (1'h1)))
            begin
              reg1068 = reg1072[(5'h11):(3'h4)];
              reg1069 = ($unsigned({{reg1056[(5'h11):(3'h7)],
                          $unsigned(reg1064)}}) ?
                  (~$signed((~&((8'hb8) ? reg1072 : reg1052)))) : (!((((8'h9c) ?
                              reg1045 : reg1059) ?
                          $unsigned(reg1069) : $signed(reg1066)) ?
                      ((~reg1035) && reg1035[(5'h10):(1'h1)]) : $signed({reg1034,
                          reg1068}))));
            end
          reg1070 = {$signed({((forvar1071 <<< reg1059) ?
                      (&reg1046) : $unsigned((8'ha0)))})};
          reg1071 = ((^~$unsigned((wire1029 ? (~|reg1073) : forvar1071))) ?
              reg1051[(4'hf):(4'hf)] : (~^(8'had)));
          reg1072 = $unsigned((+reg1073));
          for (forvar1073 = (1'h0); (forvar1073 < (2'h3)); forvar1073 = (forvar1073 + (1'h1)))
            begin
              reg1075 = (reg1032 ? reg1074[(1'h1):(1'h0)] : reg1066);
              reg1076 <= wire1054[(5'h14):(5'h13)];
              reg1077 = forvar1073[(4'he):(3'h6)];
              reg1078 = $unsigned((((8'hb8) * $unsigned($unsigned(reg1036))) >> (^~reg1063[(1'h0):(1'h0)])));
            end
        end
    end
  always
    @(posedge clk) begin
      reg1079 = ($unsigned((^$unsigned(reg1057))) ~^ ((($unsigned(reg1045) ?
              (wire1026 ? reg1049 : wire1053) : (reg1046 || wire1026)) ?
          (+reg1064[(5'h12):(3'h5)]) : $signed($unsigned((7'h4a)))) || (^$signed(reg1057[(3'h6):(3'h6)]))));
      if (reg1045)
        begin
          if ($signed($signed((~&((reg1073 >>> reg1067) ?
              (wire1053 ? wire1028 : (8'hb2)) : reg1034)))))
            begin
              reg1080 = reg1062;
              reg1081 = $unsigned($unsigned((reg1063[(3'h6):(1'h1)] ?
                  $unsigned($signed(reg1080)) : $unsigned((wire1026 ?
                      (8'hba) : reg1035)))));
              reg1082 = {(reg1064 << $unsigned((wire1030 ?
                      $signed(wire1028) : $signed(reg1039)))),
                  reg1034[(4'h9):(2'h2)]};
            end
          else
            begin
              reg1080 = ((|((reg1082 >>> (^~reg1074)) & $unsigned($unsigned(wire1026)))) ?
                  {((reg1063 >= (!wire1026)) ?
                          ((reg1082 < reg1045) < $unsigned(reg1067)) : ((^wire1028) <<< $unsigned(wire1030))),
                      reg1080} : $unsigned((~&($unsigned(reg1062) ^ (+reg1045)))));
              reg1083 <= $unsigned({$signed((~|(7'h41)))});
              reg1084 = reg1046[(2'h3):(2'h3)];
            end
          reg1085 = {$unsigned((|((wire1030 ?
                  reg1081 : reg1032) - $signed(reg1035)))),
              ((~^{(~&reg1035), reg1035[(4'hf):(4'hb)]}) ?
                  $signed(($signed(wire1029) ?
                      (~reg1039) : (reg1082 - reg1079))) : {reg1084})};
        end
      else
        begin
          for (forvar1080 = (1'h0); (forvar1080 < (1'h0)); forvar1080 = (forvar1080 + (1'h1)))
            begin
              reg1081 = {forvar1080[(2'h2):(1'h0)],
                  ((+$signed((reg1035 ? reg1062 : reg1034))) ?
                      ((8'h9c) ?
                          ((reg1073 ? (8'hb4) : reg1035) ?
                              $signed(reg1055) : (&wire1030)) : ({wire1028} || {reg1083,
                              (8'hb2)})) : (reg1041[(2'h2):(1'h1)] ?
                          (^$signed(reg1055)) : $signed((^reg1057))))};
              reg1082 = $signed({(((-wire1030) && reg1084) ^ reg1063)});
              reg1084 = $signed(reg1055);
              reg1086 <= reg1064[(1'h1):(1'h0)];
            end
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned($unsigned(reg1055)))
        begin
          if (reg1045[(5'h10):(3'h4)])
            begin
              reg1087 <= (~&{({{(8'hb9), (8'hb4)}, (reg1073 | reg1035)} ?
                      reg1034[(5'h14):(3'h4)] : reg1032[(4'hd):(3'h4)])});
              reg1088 = reg1063[(3'h4):(1'h1)];
            end
          else
            begin
              reg1088 = (reg1032 ?
                  reg1057[(3'h7):(3'h6)] : reg1039[(3'h5):(3'h5)]);
              reg1089 = reg1073;
              reg1090 <= ({(($unsigned((8'hb3)) <<< $unsigned(reg1046)) ?
                      (~|{(8'h9d)}) : (reg1074[(2'h3):(1'h1)] ^ (reg1089 && wire1053))),
                  ((7'h44) ?
                      $unsigned((wire1053 | (8'ha6))) : ({reg1057,
                          reg1083} + ((7'h40) ?
                          wire1029 : reg1041)))} <= $unsigned(((7'h46) ?
                  $unsigned({reg1039,
                      reg1088}) : ((reg1086 ^~ (8'had)) || (~&reg1049)))));
              reg1091 = (((~&reg1038[(3'h7):(1'h0)]) ?
                  (+$unsigned($unsigned(reg1052))) : $unsigned($signed(wire1030))) && $signed(reg1055));
            end
          for (forvar1092 = (1'h0); (forvar1092 < (3'h4)); forvar1092 = (forvar1092 + (1'h1)))
            begin
              reg1093 = ($unsigned(($unsigned(((8'hbb) ? (8'haa) : wire1054)) ?
                  $unsigned((reg1035 ?
                      wire1054 : reg1051)) : reg1076)) && {$unsigned($signed((~|reg1034))),
                  $unsigned(reg1052[(4'ha):(4'h8)])});
              reg1094 <= reg1052[(1'h0):(1'h0)];
              reg1095 = reg1049[(3'h4):(2'h2)];
            end
          reg1096 <= reg1036;
        end
      else
        begin
          for (forvar1087 = (1'h0); (forvar1087 < (2'h2)); forvar1087 = (forvar1087 + (1'h1)))
            begin
              reg1088 = $unsigned(({(!(8'hb2))} > (|$signed($signed(wire1026)))));
              reg1089 = $unsigned($signed(forvar1087));
            end
          if (((&(^~reg1049)) >>> reg1047))
            begin
              reg1090 <= ($signed($unsigned($signed((reg1057 <<< wire1054)))) ?
                  reg1049 : ((8'hb3) >> reg1035));
              reg1091 = ((+$signed($unsigned(((7'h4a) && reg1032)))) ?
                  reg1093 : reg1064);
            end
          else
            begin
              reg1090 <= $unsigned(reg1055[(4'h8):(3'h6)]);
            end
          reg1092 <= reg1064[(5'h13):(4'hc)];
        end
      reg1097 <= $unsigned(reg1091);
      if ((((^~reg1090[(1'h1):(1'h0)]) || $signed($signed((~reg1036)))) ?
          reg1047[(1'h1):(1'h0)] : (~&reg1095)))
        begin
          for (forvar1098 = (1'h0); (forvar1098 < (1'h0)); forvar1098 = (forvar1098 + (1'h1)))
            begin
              reg1099 <= ({{reg1076, {$unsigned(reg1086)}},
                  reg1087[(2'h2):(2'h2)]} < {((~|$unsigned(reg1064)) ?
                      {(reg1074 & reg1045)} : (&((8'h9e) ?
                          wire1029 : reg1035))),
                  (8'hb7)});
              reg1100 = $unsigned($unsigned(reg1087[(1'h1):(1'h1)]));
              reg1101 = $signed((+$signed($signed(reg1036))));
              reg1102 = (((({(8'hb0)} <<< (reg1047 || reg1038)) ?
                      $signed(((8'haf) ?
                          reg1046 : (8'ha0))) : reg1087[(2'h2):(1'h0)]) ?
                  ($signed(reg1062[(4'hd):(4'h8)]) ^ $signed({wire1027})) : wire1029[(2'h3):(2'h2)]) + $unsigned(reg1046[(3'h7):(1'h0)]));
            end
          if ({((&(reg1057 ?
                  {forvar1092, reg1046} : {reg1096})) || $signed((wire1053 ?
                  reg1063 : reg1097))),
              $unsigned($signed($unsigned((+(7'h40)))))})
            begin
              reg1103 <= (reg1067 && reg1091);
            end
          else
            begin
              reg1104 = (reg1096 ?
                  $unsigned((~^($signed(reg1092) ?
                      reg1076 : (reg1090 ?
                          (8'hb8) : (7'h48))))) : ((~|($signed(reg1095) || $unsigned(reg1095))) ?
                      (8'hb4) : (((wire1030 ? reg1051 : reg1063) > reg1083) ?
                          (^~(reg1052 ? reg1076 : wire1029)) : reg1088)));
              reg1105 <= $unsigned((~^(((+reg1073) ?
                      $unsigned(reg1102) : reg1039) ?
                  reg1083[(3'h5):(1'h1)] : (~|wire1027[(4'ha):(3'h7)]))));
            end
        end
      else
        begin
          for (forvar1098 = (1'h0); (forvar1098 < (1'h1)); forvar1098 = (forvar1098 + (1'h1)))
            begin
              reg1099 <= $signed(reg1100);
              reg1103 <= reg1057;
            end
          reg1105 <= reg1039;
          for (forvar1106 = (1'h0); (forvar1106 < (1'h1)); forvar1106 = (forvar1106 + (1'h1)))
            begin
              reg1107 = $signed((~&$unsigned((reg1086 ?
                  $unsigned(reg1089) : wire1029))));
              reg1108 = {((-forvar1106[(4'ha):(3'h6)]) >>> $signed(reg1090))};
            end
        end
      if (reg1104)
        begin
          for (forvar1109 = (1'h0); (forvar1109 < (2'h3)); forvar1109 = (forvar1109 + (1'h1)))
            begin
              reg1110 = ($unsigned((!reg1083)) ~^ reg1096[(5'h17):(2'h3)]);
              reg1111 = (reg1045 ?
                  $unsigned(reg1047) : {((forvar1098[(4'hb):(4'hb)] != $unsigned(reg1034)) ?
                          (reg1101 ?
                              reg1108[(2'h3):(2'h2)] : $signed(reg1055)) : $signed((8'ha8))),
                      $unsigned(reg1049[(1'h0):(1'h0)])});
              reg1112 = $unsigned(wire1030);
              reg1113 = $signed($signed(forvar1087));
            end
          for (forvar1114 = (1'h0); (forvar1114 < (1'h0)); forvar1114 = (forvar1114 + (1'h1)))
            begin
              reg1115 = forvar1087;
              reg1116 <= ((8'hac) ?
                  wire1030 : {reg1051[(5'h15):(4'h9)],
                      (^$unsigned($unsigned(wire1026)))});
            end
          reg1117 = (reg1093 > {reg1034});
        end
      else
        begin
          reg1109 = forvar1106;
          if ($signed(reg1035))
            begin
              reg1114 <= ({({$signed(wire1028)} >>> (~^((8'ha1) >> forvar1106)))} ?
                  ((reg1067 ?
                          ((reg1112 ? reg1074 : wire1054) ?
                              {(8'hb9)} : (~&(8'ha8))) : $unsigned($unsigned(reg1062))) ?
                      ((!$signed(forvar1106)) ?
                          reg1113[(1'h1):(1'h1)] : ((reg1102 ?
                              (8'hb0) : reg1103) & (~&forvar1114))) : reg1115) : $unsigned($signed($unsigned({forvar1106}))));
              reg1116 <= {(~|$signed(((^reg1047) ?
                      ((8'hb7) ? reg1095 : reg1076) : $unsigned((8'hb9))))),
                  ($unsigned(((reg1032 < wire1027) == (reg1105 * reg1090))) ?
                      ({{reg1064, forvar1098},
                          {reg1051}} >>> ($signed(reg1091) ?
                          $unsigned(forvar1098) : (reg1107 ?
                              (8'ha3) : reg1087))) : ((-(8'h9e)) ?
                          reg1091[(4'h8):(3'h6)] : (&reg1034)))};
              reg1118 <= forvar1109;
            end
          else
            begin
              reg1110 = reg1104[(3'h4):(1'h1)];
              reg1111 = reg1113;
              reg1114 <= ((~$unsigned(wire1027)) && {reg1100});
              reg1116 <= wire1027;
            end
        end
      reg1119 <= reg1118[(1'h1):(1'h1)];
    end
  assign wire1120 = (~((~^$unsigned((~reg1035))) ~^ (~|($unsigned(reg1073) ?
                        (8'ha9) : (reg1103 ? reg1035 : reg1074)))));
  assign wire1121 = (|$signed(reg1041));
  assign wire1122 = $signed(reg1051);
  assign wire1123 = (($signed($unsigned((wire1121 << reg1114))) ?
                            $unsigned(((wire1030 ? reg1073 : (8'haf)) ?
                                reg1074 : (reg1052 > reg1090))) : reg1064) ?
                        reg1036 : reg1034[(4'h9):(3'h6)]);
  assign wire1124 = reg1087[(3'h6):(1'h0)];
  assign wire1125 = ((^~(~(-(reg1039 == wire1054)))) ?
                        $unsigned({$unsigned(reg1063[(4'h8):(2'h3)]),
                            $unsigned($unsigned((7'h4a)))}) : ((reg1064[(4'ha):(4'h9)] ?
                            ((wire1121 ?
                                (8'h9e) : reg1046) ^~ $signed(reg1032)) : reg1096) >> wire1120[(4'h8):(3'h7)]));
  assign wire1126 = (reg1047 ?
                        ($signed(reg1116) ?
                            (+$signed($unsigned(reg1083))) : (reg1041 ?
                                reg1083[(3'h5):(3'h4)] : $unsigned((-(7'h41))))) : reg1087[(2'h3):(2'h3)]);
  always
    @(posedge clk) begin
      if ((wire1027 ? reg1036 : $unsigned((8'hb6))))
        begin
          if ($signed((wire1028 ?
              $signed(($signed(reg1039) ?
                  (^~wire1121) : {(8'ha8)})) : {$signed($unsigned(wire1027))})))
            begin
              reg1127 <= (^(-reg1114));
              reg1128 = (($unsigned(reg1094[(2'h2):(1'h0)]) ?
                  $unsigned((!(~^reg1039))) : ($unsigned($unsigned(reg1099)) || reg1038)) && ((^~{(reg1046 >>> reg1049),
                  (wire1054 < wire1121)}) + (&reg1127[(3'h7):(2'h3)])));
              reg1129 = ((reg1047 ?
                  (($signed(reg1038) ^~ (-reg1041)) & ((reg1034 ?
                      reg1096 : reg1032) | (7'h45))) : wire1027[(3'h6):(1'h1)]) | {reg1038[(3'h6):(2'h3)]});
              reg1130 = reg1099;
            end
          else
            begin
              reg1127 <= ((7'h45) ? (8'haf) : reg1105[(5'h17):(5'h12)]);
              reg1131 <= {(~&($unsigned(reg1083) ?
                      wire1027 : ((reg1073 ? wire1027 : reg1046) ?
                          $unsigned(reg1086) : $unsigned((8'ha4))))),
                  reg1041};
              reg1132 = $unsigned($unsigned({({reg1092} ~^ $unsigned((8'h9c)))}));
              reg1133 <= (reg1073 ?
                  (~{({reg1127} ?
                          $unsigned(wire1054) : $signed(reg1047))}) : (8'hb4));
            end
        end
      else
        begin
          for (forvar1127 = (1'h0); (forvar1127 < (3'h4)); forvar1127 = (forvar1127 + (1'h1)))
            begin
              reg1131 <= (reg1036[(1'h0):(1'h0)] & (wire1124[(1'h1):(1'h1)] != $signed({$signed(wire1026)})));
              reg1132 = $signed($unsigned({(wire1028 != (reg1086 * reg1096))}));
            end
          for (forvar1133 = (1'h0); (forvar1133 < (1'h1)); forvar1133 = (forvar1133 + (1'h1)))
            begin
              reg1134 = wire1053;
              reg1135 = (~&(((wire1026[(2'h3):(1'h1)] ?
                  $signed(reg1097) : (reg1096 ?
                      wire1027 : reg1062)) ~^ $signed($unsigned(reg1099))) * reg1067));
            end
          reg1136 = {reg1062};
        end
      reg1137 <= (~reg1131[(4'h9):(3'h4)]);
    end
  assign wire1138 = $unsigned((8'hb7));
  always
    @(posedge clk) begin
      for (forvar1139 = (1'h0); (forvar1139 < (3'h4)); forvar1139 = (forvar1139 + (1'h1)))
        begin
          for (forvar1140 = (1'h0); (forvar1140 < (1'h0)); forvar1140 = (forvar1140 + (1'h1)))
            begin
              reg1141 <= wire1138[(1'h0):(1'h0)];
              reg1142 = $unsigned({wire1126,
                  $signed((&(wire1122 && wire1029)))});
            end
          for (forvar1143 = (1'h0); (forvar1143 < (1'h0)); forvar1143 = (forvar1143 + (1'h1)))
            begin
              reg1144 <= {(~(~(reg1067[(3'h6):(1'h1)] >= (reg1083 ?
                      reg1051 : (8'hab))))),
                  $unsigned((8'hb1))};
            end
          if (wire1124)
            begin
              reg1145 = (reg1141 <= (wire1121[(3'h6):(3'h5)] || ($signed($unsigned(wire1122)) >> reg1133[(4'hb):(2'h3)])));
            end
          else
            begin
              reg1145 = reg1057[(3'h7):(3'h7)];
              reg1146 <= (8'hae);
              reg1147 = {(8'hab), wire1026[(2'h3):(1'h1)]};
            end
          for (forvar1148 = (1'h0); (forvar1148 < (2'h2)); forvar1148 = (forvar1148 + (1'h1)))
            begin
              reg1149 = ($signed($signed(reg1038)) ?
                  $unsigned(({((8'hb7) ? reg1133 : reg1118),
                          {reg1076, reg1114}} ?
                      ((reg1133 ? wire1138 : reg1035) >= {reg1097,
                          wire1030}) : $unsigned(reg1142))) : $signed($unsigned(reg1105[(4'h8):(3'h6)])));
              reg1150 <= ($signed($signed(reg1092)) >>> ((reg1092 ?
                      $unsigned(reg1067) : reg1103[(5'h16):(4'h8)]) ?
                  (reg1047 && reg1034) : $signed(wire1030[(1'h0):(1'h0)])));
              reg1151 = ($unsigned((reg1064[(3'h7):(3'h7)] ?
                  $unsigned((wire1124 <= wire1123)) : (&$signed(reg1083)))) < ($unsigned($unsigned((-reg1046))) + $signed(((reg1067 ?
                  reg1062 : (8'hb3)) >= $unsigned(wire1028)))));
              reg1152 <= wire1028[(1'h1):(1'h0)];
              reg1153 <= $unsigned(reg1052);
            end
          for (forvar1154 = (1'h0); (forvar1154 < (3'h4)); forvar1154 = (forvar1154 + (1'h1)))
            begin
              reg1155 = (~^((8'ha8) <<< ($signed((wire1122 || reg1149)) << (&$signed(reg1076)))));
              reg1156 = $signed(($unsigned($unsigned($signed(reg1038))) << {{(wire1138 ?
                          reg1152 : (7'h46)),
                      (~&reg1052)}}));
              reg1157 = $signed($unsigned(((^~{reg1133,
                  wire1028}) >= $unsigned($signed((8'hbf))))));
              reg1158 = (^~(reg1034[(2'h2):(1'h1)] || $unsigned($unsigned($unsigned(wire1125)))));
            end
        end
      reg1159 = ((^$signed((~&{reg1067, (7'h42)}))) ?
          $signed(reg1141[(1'h1):(1'h0)]) : reg1046);
      for (forvar1160 = (1'h0); (forvar1160 < (2'h2)); forvar1160 = (forvar1160 + (1'h1)))
        begin
          reg1161 <= (~&$unsigned(reg1158));
          if (({reg1062} ?
              ((7'h43) | (&$unsigned((reg1133 ?
                  reg1035 : reg1145)))) : (7'h41)))
            begin
              reg1162 = ((reg1131 ?
                  ((&$signed(reg1046)) < $signed((reg1032 ^~ reg1131))) : $signed(reg1151[(4'hb):(2'h3)])) >>> $unsigned(((8'haa) | $unsigned(wire1124))));
              reg1163 <= (reg1064[(5'h12):(5'h11)] > {(($unsigned(reg1083) ?
                      $signed(reg1127) : wire1054[(3'h4):(1'h1)]) + $signed((reg1045 ?
                      reg1105 : reg1052))),
                  reg1144[(2'h3):(2'h3)]});
              reg1164 <= $unsigned($unsigned(($unsigned({wire1120, reg1052}) ?
                  (-$unsigned(reg1161)) : {$unsigned(reg1163)})));
            end
          else
            begin
              reg1162 = {$signed($signed(reg1164)),
                  $unsigned($unsigned(($unsigned(reg1036) << (reg1119 & reg1051))))};
            end
          reg1165 = (reg1087 ?
              reg1145 : (reg1164[(4'hf):(4'hf)] ?
                  (^~$unsigned(reg1147[(5'h11):(4'ha)])) : $unsigned((7'h42))));
        end
      reg1166 <= $unsigned((-($unsigned(reg1094[(1'h1):(1'h0)]) ?
          $unsigned(wire1123) : ($signed((8'hbb)) <= (~|reg1074)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module863
#(parameter param993 = ((~{(((8'hae) > (7'h4a)) ~^ ((7'h4a) << (8'hb2))), (((8'hbc) ? (8'ha1) : (7'h43)) >= (~|(8'h9f)))}) ? (((((7'h44) ? (8'hb9) : (7'h48)) >> ((8'h9f) > (8'hb9))) ? (((8'hbc) || (8'ha5)) && (&(8'hab))) : {((8'haa) <<< (8'ha5)), ((8'hbc) > (7'h45))}) || (8'ha0)) : (^(~|((8'hbf) == ((8'ha0) + (8'ha4)))))))
(y, clk, wire867, wire866, wire865, wire864);
  output wire [(32'h6ef):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'h8):(1'h0)] wire867;
  input wire signed [(4'hd):(1'h0)] wire866;
  input wire [(5'h16):(1'h0)] wire865;
  input wire signed [(5'h11):(1'h0)] wire864;
  wire [(3'h6):(1'h0)] wire914;
  wire signed [(2'h3):(1'h0)] wire913;
  wire signed [(3'h4):(1'h0)] wire912;
  wire signed [(3'h4):(1'h0)] wire901;
  wire signed [(5'h17):(1'h0)] wire900;
  wire [(4'he):(1'h0)] wire870;
  wire [(3'h6):(1'h0)] wire869;
  wire [(5'h13):(1'h0)] wire868;
  reg signed [(4'hc):(1'h0)] reg991 = (1'h0);
  reg [(4'ha):(1'h0)] reg990 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg987 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg985 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg984 = (1'h0);
  reg [(5'h10):(1'h0)] reg983 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg982 = (1'h0);
  reg signed [(4'he):(1'h0)] reg980 = (1'h0);
  reg [(5'h17):(1'h0)] reg977 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg975 = (1'h0);
  reg [(3'h4):(1'h0)] reg974 = (1'h0);
  reg [(5'h17):(1'h0)] reg970 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg969 = (1'h0);
  reg [(4'hd):(1'h0)] reg967 = (1'h0);
  reg signed [(4'he):(1'h0)] reg964 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg963 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg962 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg961 = (1'h0);
  reg [(4'hf):(1'h0)] reg959 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg956 = (1'h0);
  reg [(5'h17):(1'h0)] reg955 = (1'h0);
  reg [(5'h16):(1'h0)] reg954 = (1'h0);
  reg [(3'h5):(1'h0)] reg950 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg948 = (1'h0);
  reg [(3'h7):(1'h0)] reg946 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg945 = (1'h0);
  reg [(5'h17):(1'h0)] reg944 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg943 = (1'h0);
  reg [(5'h11):(1'h0)] reg941 = (1'h0);
  reg [(5'h18):(1'h0)] reg940 = (1'h0);
  reg [(4'hd):(1'h0)] reg939 = (1'h0);
  reg [(5'h13):(1'h0)] reg936 = (1'h0);
  reg [(4'hf):(1'h0)] reg932 = (1'h0);
  reg [(5'h17):(1'h0)] reg933 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg930 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg928 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg923 = (1'h0);
  reg [(2'h3):(1'h0)] reg922 = (1'h0);
  reg [(5'h14):(1'h0)] reg919 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg918 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg917 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg911 = (1'h0);
  reg [(3'h4):(1'h0)] reg910 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg908 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg905 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg904 = (1'h0);
  reg [(5'h15):(1'h0)] reg902 = (1'h0);
  reg [(4'h8):(1'h0)] reg891 = (1'h0);
  reg [(5'h12):(1'h0)] reg897 = (1'h0);
  reg signed [(4'he):(1'h0)] reg895 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg890 = (1'h0);
  reg [(5'h10):(1'h0)] reg888 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg887 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg883 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg879 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg877 = (1'h0);
  reg [(5'h14):(1'h0)] reg876 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg874 = (1'h0);
  reg [(3'h4):(1'h0)] reg873 = (1'h0);
  reg [(4'he):(1'h0)] reg992 = (1'h0);
  reg [(4'hb):(1'h0)] reg989 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg988 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg986 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar982 = (1'h0);
  reg [(5'h13):(1'h0)] reg978 = (1'h0);
  reg [(5'h17):(1'h0)] forvar977 = (1'h0);
  reg [(4'h9):(1'h0)] reg981 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg979 = (1'h0);
  reg [(5'h13):(1'h0)] forvar978 = (1'h0);
  reg [(4'hd):(1'h0)] reg976 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg973 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg972 = (1'h0);
  reg [(4'hd):(1'h0)] reg971 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg968 = (1'h0);
  reg [(5'h16):(1'h0)] reg966 = (1'h0);
  reg [(5'h13):(1'h0)] reg965 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg960 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg957 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar954 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg958 = (1'h0);
  reg [(4'hf):(1'h0)] forvar957 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg953 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar952 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg951 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg949 = (1'h0);
  reg [(4'hf):(1'h0)] reg947 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg942 = (1'h0);
  reg [(4'h9):(1'h0)] reg938 = (1'h0);
  reg [(2'h3):(1'h0)] forvar937 = (1'h0);
  reg [(2'h2):(1'h0)] reg935 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar931 = (1'h0);
  reg [(5'h16):(1'h0)] reg934 = (1'h0);
  reg [(4'h9):(1'h0)] forvar932 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg931 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg929 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg927 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg926 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg925 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg924 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg915 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg921 = (1'h0);
  reg [(5'h11):(1'h0)] reg920 = (1'h0);
  reg [(2'h3):(1'h0)] reg916 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar915 = (1'h0);
  reg [(5'h16):(1'h0)] reg909 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg907 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg906 = (1'h0);
  reg [(4'hc):(1'h0)] reg903 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg899 = (1'h0);
  reg [(5'h18):(1'h0)] reg898 = (1'h0);
  reg [(3'h5):(1'h0)] reg896 = (1'h0);
  reg [(3'h6):(1'h0)] forvar894 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg893 = (1'h0);
  reg [(4'hd):(1'h0)] reg892 = (1'h0);
  reg [(2'h3):(1'h0)] forvar891 = (1'h0);
  reg [(5'h17):(1'h0)] reg889 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg886 = (1'h0);
  reg [(5'h15):(1'h0)] reg885 = (1'h0);
  reg [(3'h7):(1'h0)] reg884 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg882 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg881 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar876 = (1'h0);
  reg [(5'h17):(1'h0)] reg880 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg878 = (1'h0);
  reg [(5'h17):(1'h0)] reg875 = (1'h0);
  reg [(5'h11):(1'h0)] reg872 = (1'h0);
  reg [(4'hc):(1'h0)] reg871 = (1'h0);
  assign y = {wire914,
                 wire913,
                 wire912,
                 wire901,
                 wire900,
                 wire870,
                 wire869,
                 wire868,
                 reg991,
                 reg990,
                 reg987,
                 reg985,
                 reg984,
                 reg983,
                 reg982,
                 reg980,
                 reg977,
                 reg975,
                 reg974,
                 reg970,
                 reg969,
                 reg967,
                 reg964,
                 reg963,
                 reg962,
                 reg961,
                 reg959,
                 reg956,
                 reg955,
                 reg954,
                 reg950,
                 reg948,
                 reg946,
                 reg945,
                 reg944,
                 reg943,
                 reg941,
                 reg940,
                 reg939,
                 reg936,
                 reg932,
                 reg933,
                 reg930,
                 reg928,
                 reg923,
                 reg922,
                 reg919,
                 reg918,
                 reg917,
                 reg911,
                 reg910,
                 reg908,
                 reg905,
                 reg904,
                 reg902,
                 reg891,
                 reg897,
                 reg895,
                 reg890,
                 reg888,
                 reg887,
                 reg883,
                 reg879,
                 reg877,
                 reg876,
                 reg874,
                 reg873,
                 reg992,
                 reg989,
                 reg988,
                 reg986,
                 forvar982,
                 reg978,
                 forvar977,
                 reg981,
                 reg979,
                 forvar978,
                 reg976,
                 reg973,
                 reg972,
                 reg971,
                 reg968,
                 reg966,
                 reg965,
                 reg960,
                 reg957,
                 forvar954,
                 reg958,
                 forvar957,
                 reg953,
                 forvar952,
                 reg951,
                 reg949,
                 reg947,
                 reg942,
                 reg938,
                 forvar937,
                 reg935,
                 forvar931,
                 reg934,
                 forvar932,
                 reg931,
                 reg929,
                 reg927,
                 reg926,
                 reg925,
                 reg924,
                 reg915,
                 reg921,
                 reg920,
                 reg916,
                 forvar915,
                 reg909,
                 reg907,
                 reg906,
                 reg903,
                 reg899,
                 reg898,
                 reg896,
                 forvar894,
                 reg893,
                 reg892,
                 forvar891,
                 reg889,
                 reg886,
                 reg885,
                 reg884,
                 reg882,
                 reg881,
                 forvar876,
                 reg880,
                 reg878,
                 reg875,
                 reg872,
                 reg871,
                 (1'h0)};
  assign wire868 = (({$signed($signed(wire864))} ?
                       $unsigned((8'ha4)) : $signed($unsigned($signed(wire866)))) ^~ (8'ha4));
  assign wire869 = wire868;
  assign wire870 = (^~((wire867[(3'h5):(2'h2)] ?
                       (wire868[(3'h6):(3'h6)] ?
                           (+(8'hac)) : $unsigned((8'ha8))) : wire864) > (8'hb1)));
  always
    @(posedge clk) begin
      reg871 = $unsigned((wire868[(4'hd):(3'h5)] ?
          wire869[(2'h3):(1'h1)] : $unsigned(wire868)));
      reg872 = $signed(wire865);
    end
  always
    @(posedge clk) begin
      if (($unsigned($unsigned((wire867[(4'h8):(3'h6)] ?
          wire868 : {(7'h48)}))) != {wire866[(1'h1):(1'h0)]}))
        begin
          if (wire870)
            begin
              reg873 <= (wire870 ? wire869 : wire869);
              reg874 <= (!$unsigned($unsigned($signed(reg873[(1'h1):(1'h0)]))));
            end
          else
            begin
              reg875 = ((reg873 * (reg873 ?
                      (^~(reg874 ? wire869 : wire870)) : (^~(^reg874)))) ?
                  (^reg874) : $signed(((wire865[(4'hf):(3'h7)] ?
                          (wire868 <<< wire868) : (wire869 != (8'ha7))) ?
                      wire865[(4'hc):(4'hc)] : (^~wire867[(1'h1):(1'h0)]))));
              reg876 <= $signed($unsigned((((wire870 != wire867) ?
                      (&wire866) : (^wire864)) ?
                  $unsigned(reg875) : reg874)));
              reg877 <= ((wire870 ?
                      ($unsigned({reg874,
                          wire865}) || wire867[(3'h7):(3'h5)]) : (wire867[(3'h4):(1'h1)] + (((8'had) ?
                              wire867 : reg876) ?
                          $signed((8'ha8)) : (wire870 ? reg875 : reg875)))) ?
                  (+reg874) : (8'h9c));
              reg878 = $signed($unsigned({reg875[(4'hd):(3'h6)],
                  $unsigned($signed(reg875))}));
            end
          if ({{$signed(($unsigned(reg877) ?
                      (wire865 - wire869) : reg875[(4'hc):(4'ha)])),
                  {((&(8'hb9)) != (8'h9d))}},
              $signed(wire866[(4'h9):(2'h3)])})
            begin
              reg879 <= wire870;
            end
          else
            begin
              reg880 = {{wire867, wire869},
                  (reg875 ?
                      (^~{(reg873 <= wire864)}) : (reg874[(1'h1):(1'h0)] ~^ (reg878 ?
                          reg878 : $unsigned(reg878))))};
            end
        end
      else
        begin
          reg875 = (~|(!(8'hbb)));
          for (forvar876 = (1'h0); (forvar876 < (2'h2)); forvar876 = (forvar876 + (1'h1)))
            begin
              reg877 <= ((~|reg879[(4'h8):(3'h5)]) ?
                  ((~^$signed(((8'hbb) <= reg876))) ^~ reg877) : $signed($unsigned((8'hbb))));
              reg878 = (7'h4a);
            end
          reg880 = (({$unsigned($unsigned((8'hbf)))} ? wire864 : wire868) ?
              ({(((8'h9c) ? wire865 : reg875) ? {reg874} : reg876),
                  (|((8'hac) * wire870))} <= (~&{$signed((8'hb1))})) : reg874[(3'h4):(2'h2)]);
          if ($unsigned((^~{(+$unsigned(forvar876)),
              (&(wire868 ? reg875 : reg880))})))
            begin
              reg881 = {(+reg876)};
              reg882 = ($signed($unsigned($unsigned((+reg881)))) == ((-((wire866 ^ (8'hb4)) ?
                  wire865[(5'h16):(5'h13)] : (8'hab))) >= wire868));
              reg883 <= $signed(reg875);
            end
          else
            begin
              reg881 = $unsigned(wire864[(4'hd):(4'hd)]);
              reg882 = wire869[(3'h5):(3'h5)];
              reg884 = (~^((wire870 ?
                      $unsigned(reg883[(2'h2):(2'h2)]) : {(~^reg877)}) ?
                  (~$signed(reg880[(1'h1):(1'h1)])) : $unsigned((7'h48))));
              reg885 = wire868[(4'h9):(4'h8)];
              reg886 = $signed(($signed($unsigned(reg884)) ? reg885 : wire869));
            end
          reg887 <= $signed($signed(reg880[(1'h1):(1'h1)]));
        end
      reg888 <= $signed((|$signed(($signed(wire869) + wire864[(4'he):(4'ha)]))));
      reg889 = ($unsigned(reg879) & {$unsigned((reg880[(1'h0):(1'h0)] < $unsigned(wire868))),
          (-$signed((!wire865)))});
      reg890 <= (reg882[(1'h1):(1'h0)] ?
          (reg879[(4'hd):(2'h3)] ?
              {$unsigned(reg873)} : (~|$signed(wire864))) : $signed(reg889));
      if ((|(+{((forvar876 <= wire867) ?
              $unsigned((8'had)) : $unsigned(reg877))})))
        begin
          for (forvar891 = (1'h0); (forvar891 < (1'h0)); forvar891 = (forvar891 + (1'h1)))
            begin
              reg892 = reg885[(1'h0):(1'h0)];
            end
          reg893 = (!$signed(((+wire868[(3'h5):(3'h5)]) ?
              reg875[(4'h8):(3'h4)] : (~(7'h41)))));
          for (forvar894 = (1'h0); (forvar894 < (3'h4)); forvar894 = (forvar894 + (1'h1)))
            begin
              reg895 <= $signed((~^wire866[(4'hc):(4'h8)]));
              reg896 = $unsigned(((reg875[(4'h8):(1'h1)] ?
                  (((8'hae) ? reg880 : reg876) ?
                      $unsigned(reg873) : (reg893 | reg882)) : {reg893[(3'h7):(2'h3)]}) == (((|reg880) ?
                      (reg875 ? reg878 : reg879) : wire864[(3'h7):(3'h5)]) ?
                  reg885 : {{wire867}, forvar894[(1'h0):(1'h0)]})));
              reg897 <= (^($signed((8'hae)) ?
                  $signed(reg886) : $unsigned($unsigned($signed((7'h45))))));
              reg898 = $signed(((~reg883[(1'h1):(1'h1)]) == reg885[(4'hd):(1'h1)]));
              reg899 = $unsigned((reg889 >>> forvar891[(2'h2):(1'h1)]));
            end
        end
      else
        begin
          reg891 <= ($unsigned(($signed((reg875 ?
                  reg874 : reg873)) ~^ {$unsigned((8'hb8))})) ?
              {($signed((forvar891 ? wire864 : reg879)) ?
                      {(~&(8'hbf))} : reg884[(3'h4):(2'h3)])} : reg895);
        end
    end
  assign wire900 = $unsigned(reg895);
  assign wire901 = reg874;
  always
    @(posedge clk) begin
      if ((&wire900[(5'h15):(3'h5)]))
        begin
          reg902 <= ($unsigned(wire868) ?
              (&$unsigned((-$unsigned(wire900)))) : ($signed((7'h42)) ?
                  ({{wire866}} ?
                      $unsigned((~(7'h48))) : (8'hb0)) : ($unsigned((wire901 ?
                      reg877 : (8'hb9))) + wire901[(2'h3):(1'h0)])));
        end
      else
        begin
          if ((-wire900))
            begin
              reg903 = {reg876[(3'h6):(1'h0)]};
              reg904 <= (~|wire866[(3'h6):(2'h3)]);
              reg905 <= $unsigned({(^~(^$signed(reg877)))});
            end
          else
            begin
              reg903 = $unsigned($unsigned(wire868));
            end
          if (wire867)
            begin
              reg906 = (|(8'hae));
              reg907 = wire869;
              reg908 <= ((^~(($signed(wire870) || (~^wire866)) ?
                      ($signed(reg890) ?
                          $unsigned(wire866) : $signed(reg907)) : (~(reg904 >> reg902)))) ?
                  ((~&$unsigned($unsigned((8'hb7)))) | $signed((reg897 ?
                      (^reg897) : (reg877 ?
                          reg874 : (7'h41))))) : ($unsigned({wire901[(2'h2):(1'h0)]}) ?
                      (^~wire900[(5'h11):(5'h11)]) : $signed(reg879)));
              reg909 = ($unsigned((8'hae)) == wire901[(3'h4):(1'h0)]);
              reg910 <= reg891;
            end
          else
            begin
              reg908 <= reg897;
              reg910 <= $signed(($unsigned(reg903[(4'hc):(4'hc)]) == ($unsigned({wire866,
                  reg904}) >= {(wire869 >> (7'h42))})));
            end
          reg911 <= ((-($unsigned(reg883) ?
              $signed($unsigned(wire865)) : (~&{reg879,
                  wire866}))) * $signed({($signed((8'h9c)) != $unsigned(reg903))}));
        end
    end
  assign wire912 = (~^$signed($signed($signed((!(8'hbe))))));
  assign wire913 = wire901;
  assign wire914 = $signed((reg895[(2'h3):(1'h1)] ?
                       (^(8'hb2)) : (!$unsigned($signed(reg891)))));
  always
    @(posedge clk) begin
      if (reg897[(5'h12):(4'hc)])
        begin
          for (forvar915 = (1'h0); (forvar915 < (2'h3)); forvar915 = (forvar915 + (1'h1)))
            begin
              reg916 = $signed(reg877[(4'he):(1'h1)]);
            end
          if ($signed(forvar915[(3'h7):(2'h2)]))
            begin
              reg917 <= $signed($signed($unsigned(wire900[(3'h4):(3'h4)])));
              reg918 <= {$signed((&($unsigned(wire914) ?
                      $signed(reg904) : $unsigned((8'had)))))};
              reg919 <= (~^(^~$unsigned((8'hb5))));
              reg920 = (((~^{$unsigned((8'hbd))}) >> ($signed(reg918) + reg890[(4'h8):(4'h8)])) ?
                  wire866 : ((-(8'hb4)) ?
                      ((~{reg895}) ?
                          $unsigned(reg917[(1'h1):(1'h1)]) : (forvar915 ?
                              {reg910,
                                  wire901} : $signed(wire901))) : reg890[(1'h1):(1'h0)]));
            end
          else
            begin
              reg917 <= (|(~^$signed(wire868[(4'hb):(3'h7)])));
              reg918 <= $signed($unsigned({(~^forvar915)}));
            end
          if ((!(($signed(((8'ha8) ? reg911 : (8'hbb))) ?
                  $signed((reg876 * wire865)) : {$unsigned(reg920)}) ?
              wire869[(1'h0):(1'h0)] : $signed($signed((wire865 << reg888))))))
            begin
              reg921 = $signed((-$unsigned($signed($signed(reg891)))));
            end
          else
            begin
              reg922 <= $unsigned(reg873);
              reg923 <= ($unsigned(((reg891 ?
                  (!reg918) : (reg883 || reg908)) ^~ $signed((wire867 ?
                  wire866 : reg904)))) == wire865);
            end
        end
      else
        begin
          if (reg887[(4'hc):(2'h2)])
            begin
              reg915 = {wire869,
                  (~(($signed(forvar915) ^ (reg890 > reg897)) || (~^wire913[(2'h3):(1'h0)])))};
              reg916 = reg890;
              reg917 <= (8'ha9);
              reg918 <= reg917[(2'h2):(1'h1)];
              reg919 <= ($signed($signed(reg890)) | $unsigned((^~{$signed(wire900)})));
            end
          else
            begin
              reg915 = reg879;
              reg917 <= {reg891[(4'h8):(2'h2)]};
              reg920 = reg890;
              reg921 = (^(7'h49));
              reg922 <= {((~&$unsigned((wire912 ? reg921 : reg922))) ?
                      {reg883[(1'h0):(1'h0)],
                          reg908[(4'h9):(3'h5)]} : (|(~^(^wire869))))};
            end
          if ((((reg917 ? (reg902 < (reg911 ^ wire868)) : reg923) ?
                  (&wire866) : (wire865 == $unsigned(((8'hae) ?
                      (8'ha4) : wire913)))) ?
              {reg915,
                  $signed($signed(reg904[(4'hb):(2'h3)]))} : $signed($unsigned(($unsigned(wire912) + (|reg879))))))
            begin
              reg924 = wire870[(3'h6):(2'h2)];
              reg925 = wire900[(1'h1):(1'h0)];
              reg926 = reg883[(1'h1):(1'h1)];
              reg927 = (~^(~wire913));
              reg928 <= reg927;
            end
          else
            begin
              reg924 = {(($unsigned($signed(reg873)) ?
                          ((reg905 > (7'h47)) ?
                              (-reg917) : (wire914 ?
                                  (7'h44) : wire870)) : ((reg883 ?
                              reg897 : reg921) != $signed(reg911))) ?
                      (reg915 ?
                          $unsigned($signed((8'ha4))) : (&wire865)) : $unsigned($signed($signed(reg902))))};
              reg928 <= ($signed(reg905[(3'h5):(2'h3)]) ^~ {reg879});
            end
          reg929 = ($signed((reg918 ? wire866[(4'hb):(1'h1)] : reg927)) ?
              (7'h48) : ((reg895[(3'h5):(3'h4)] ?
                  {reg928[(3'h4):(2'h3)],
                      $signed(reg917)} : $unsigned((8'hae))) >>> (wire868 ~^ (8'hbd))));
          reg930 <= (~|{reg922[(2'h3):(2'h3)]});
        end
      if (reg925)
        begin
          reg931 = $signed(($unsigned(($signed(reg926) ~^ (!(8'h9e)))) || ({(^~reg876)} & (reg888 + $signed(wire864)))));
          for (forvar932 = (1'h0); (forvar932 < (3'h4)); forvar932 = (forvar932 + (1'h1)))
            begin
              reg933 <= $signed(reg923[(4'ha):(4'h8)]);
              reg934 = reg924[(2'h3):(1'h1)];
            end
        end
      else
        begin
          for (forvar931 = (1'h0); (forvar931 < (3'h4)); forvar931 = (forvar931 + (1'h1)))
            begin
              reg932 <= (^reg916[(2'h2):(2'h2)]);
              reg934 = (~&$signed(($unsigned($signed(forvar915)) ?
                  $signed($unsigned(wire870)) : ((reg916 ? reg895 : wire912) ?
                      (-(8'ha0)) : $signed(reg918)))));
              reg935 = wire865;
              reg936 <= reg873[(1'h1):(1'h0)];
            end
          for (forvar937 = (1'h0); (forvar937 < (2'h2)); forvar937 = (forvar937 + (1'h1)))
            begin
              reg938 = reg917;
              reg939 <= (^~((wire914 ?
                      $unsigned(((8'hae) ?
                          reg910 : reg924)) : $unsigned(reg927)) ?
                  $signed((|(~reg887))) : $signed(reg910[(3'h4):(3'h4)])));
              reg940 <= $unsigned($signed($unsigned(((reg876 == (7'h42)) & (reg935 ?
                  reg911 : wire901)))));
              reg941 <= ($signed((reg911 <<< $unsigned($unsigned(forvar915)))) ?
                  {$unsigned(reg908[(3'h4):(2'h3)]),
                      $unsigned($unsigned((reg888 || reg917)))} : {((^~(!reg895)) > reg938)});
            end
          if ({reg876, (7'h41)})
            begin
              reg942 = ((wire868 == ((~^(reg921 ? reg897 : reg936)) ?
                      reg938 : ((8'hb9) == (~&forvar932)))) ?
                  $unsigned((reg873 || (^(forvar932 & (7'h49))))) : $unsigned((((forvar937 + (7'h42)) ?
                          (!reg915) : $signed((8'hb4))) ?
                      (8'h9c) : (+(-(8'ha3))))));
              reg943 <= ({$signed((^~(~^(8'h9e)))), forvar932[(4'h9):(2'h3)]} ?
                  reg873[(2'h2):(2'h2)] : $unsigned(reg941[(5'h11):(4'hf)]));
              reg944 <= wire865[(2'h3):(2'h2)];
              reg945 <= (reg926[(1'h0):(1'h0)] >>> reg939);
              reg946 <= $signed((^~$signed(wire912[(1'h1):(1'h0)])));
            end
          else
            begin
              reg942 = ({reg911} ?
                  ((~(~&reg911[(4'h9):(4'h9)])) != $signed(({reg931, reg873} ?
                      {reg928} : wire914))) : ((8'hb6) >= ($unsigned((reg929 <= reg915)) ~^ (~^{wire901,
                      reg928}))));
              reg947 = $unsigned((^(^reg929[(1'h0):(1'h0)])));
              reg948 <= (forvar937 ?
                  (((+$signed(reg919)) >= (&(8'ha8))) ?
                      reg897 : (+(!reg939))) : wire869[(2'h2):(1'h0)]);
              reg949 = reg905;
            end
          reg950 <= reg926[(4'h8):(2'h3)];
        end
      reg951 = $signed($unsigned(reg890[(3'h6):(2'h2)]));
      for (forvar952 = (1'h0); (forvar952 < (3'h4)); forvar952 = (forvar952 + (1'h1)))
        begin
          reg953 = (^~($unsigned((|reg874[(2'h3):(1'h0)])) >> reg934[(5'h12):(3'h6)]));
        end
    end
  always
    @(posedge clk) begin
      if (reg887[(1'h1):(1'h1)])
        begin
          reg954 <= (7'h46);
          if ((reg945 ?
              $signed((~&(-{reg910}))) : (~$signed(($signed(reg945) ?
                  {reg874, reg923} : $signed(reg883))))))
            begin
              reg955 <= $unsigned(reg941);
            end
          else
            begin
              reg955 <= $unsigned($unsigned(((8'hbe) ?
                  (&$signed(reg950)) : wire869[(3'h4):(2'h3)])));
              reg956 <= $signed((8'hb3));
            end
          for (forvar957 = (1'h0); (forvar957 < (1'h1)); forvar957 = (forvar957 + (1'h1)))
            begin
              reg958 = $unsigned(reg877);
            end
        end
      else
        begin
          for (forvar954 = (1'h0); (forvar954 < (3'h4)); forvar954 = (forvar954 + (1'h1)))
            begin
              reg957 = reg922[(2'h3):(2'h3)];
              reg959 <= $unsigned(reg874[(3'h6):(3'h6)]);
              reg960 = $unsigned(reg959[(4'hc):(4'hb)]);
            end
          reg961 <= (^((($unsigned(wire900) < {wire870, (8'hb4)}) ?
                  ((~reg950) ? reg919 : (+(8'hbf))) : wire864[(3'h7):(1'h0)]) ?
              (~^$unsigned($signed(reg940))) : reg941));
          reg962 <= forvar957[(1'h1):(1'h1)];
          reg963 <= reg908;
        end
      reg964 <= $signed($unsigned(reg883));
      if ($signed(((~^reg961[(2'h2):(2'h2)]) ?
          (((reg955 ? reg933 : reg922) ?
                  $signed(reg891) : reg904[(5'h15):(3'h5)]) ?
              (7'h47) : reg943[(1'h0):(1'h0)]) : (wire912 - (reg962 ?
              {reg956} : ((8'hab) ? (8'hb5) : reg944))))))
        begin
          reg965 = (&((reg961 >> (reg918 >> (^reg943))) << $signed($signed($unsigned(reg940)))));
          reg966 = {reg897};
        end
      else
        begin
          if ((((~&wire870[(3'h7):(1'h0)]) ?
              (~&(|(reg887 ?
                  reg965 : reg895))) : $signed(reg888)) == (+reg946[(3'h6):(2'h3)])))
            begin
              reg965 = {((((~^reg873) & (reg928 >= (8'hb4))) ~^ ($signed(reg941) > $unsigned((8'h9c)))) > (^~((^(8'hb2)) <<< wire865[(4'ha):(3'h4)]))),
                  $unsigned(reg940)};
            end
          else
            begin
              reg965 = $signed(((reg895 ?
                  ((reg933 != reg940) ?
                      reg918[(4'h8):(1'h0)] : $signed(reg946)) : reg965) != (reg958[(4'hf):(4'hd)] ?
                  $unsigned(reg941) : (wire900 ?
                      reg963[(4'ha):(3'h6)] : $unsigned(wire867)))));
              reg967 <= (reg963 ? reg930 : $unsigned((7'h49)));
              reg968 = (reg877[(2'h3):(1'h1)] <= ($unsigned({(reg902 <<< reg958),
                      (8'ha4)}) ?
                  ($unsigned(((8'hab) >> wire869)) ?
                      $signed($signed((8'hbc))) : $signed((reg965 ?
                          (7'h49) : (8'h9d)))) : ($signed($unsigned(wire901)) >> $signed(reg922))));
              reg969 <= reg887;
            end
          if ((~(~^reg928)))
            begin
              reg970 <= $signed(((reg963 ?
                      ((~|reg946) ?
                          {(8'ha1),
                              reg879} : $signed(reg954)) : reg873[(2'h2):(1'h1)]) ?
                  (^$unsigned(reg930)) : (^reg945)));
            end
          else
            begin
              reg971 = (~&$unsigned(reg959));
            end
          reg972 = $unsigned($unsigned($signed(reg964)));
        end
      reg973 = reg971;
    end
  always
    @(posedge clk) begin
      reg974 <= ((^~(~&$unsigned((~&reg955)))) * reg930[(4'h8):(3'h6)]);
      reg975 <= ((^~(reg940 ?
          $unsigned({reg888, reg940}) : wire868)) | wire869[(3'h4):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg976 = (({(reg890[(3'h5):(2'h2)] >= reg962),
          $signed(reg904[(1'h0):(1'h0)])} + {reg888[(3'h7):(1'h1)]}) >> reg946);
      if ($unsigned((wire870 ? $signed($signed(reg905)) : (8'hb3))))
        begin
          reg977 <= reg918[(2'h2):(1'h1)];
          for (forvar978 = (1'h0); (forvar978 < (2'h2)); forvar978 = (forvar978 + (1'h1)))
            begin
              reg979 = reg976[(3'h5):(2'h2)];
            end
          reg980 <= $signed($unsigned((7'h45)));
          if (reg876)
            begin
              reg981 = $unsigned((+$signed((reg955[(4'he):(4'ha)] & {reg911,
                  reg940}))));
              reg982 <= $unsigned(((((~^reg933) ?
                      $unsigned(wire901) : $signed(reg923)) ?
                  (7'h48) : ($signed(reg954) ?
                      {reg905} : $signed(reg917))) * reg961[(4'hc):(1'h0)]));
              reg983 <= reg941[(4'hd):(3'h7)];
              reg984 <= ($signed($signed((reg944[(5'h17):(2'h2)] - (reg879 ?
                  reg908 : reg979)))) ^ ($signed({{reg874, reg974}, {reg940}}) ?
                  (reg891[(1'h1):(1'h1)] >= $unsigned(reg967[(2'h2):(2'h2)])) : $signed((^(wire914 ?
                      reg930 : wire866)))));
              reg985 <= $signed($signed((8'h9d)));
            end
          else
            begin
              reg981 = reg933[(1'h0):(1'h0)];
            end
        end
      else
        begin
          for (forvar977 = (1'h0); (forvar977 < (1'h0)); forvar977 = (forvar977 + (1'h1)))
            begin
              reg978 = reg897;
              reg979 = wire864;
              reg980 <= wire900;
              reg981 = wire864;
            end
          for (forvar982 = (1'h0); (forvar982 < (2'h3)); forvar982 = (forvar982 + (1'h1)))
            begin
              reg983 <= forvar977;
              reg984 <= reg917[(4'hb):(1'h1)];
            end
          if ($unsigned($unsigned(((&wire864[(4'h8):(3'h5)]) > $signed((reg969 >> reg930))))))
            begin
              reg985 <= ((|({$signed(reg959), $signed(wire864)} ?
                  (((8'hba) != reg923) ?
                      {reg946, reg985} : $signed(reg976)) : ((~(7'h44)) ?
                      {wire914,
                          reg911} : (^~reg917)))) >> $unsigned(({(!reg873)} ?
                  reg890[(3'h5):(3'h5)] : (~|$signed(wire914)))));
              reg986 = reg890;
              reg987 <= (~&reg877[(4'hf):(3'h7)]);
              reg988 = $unsigned(forvar982);
              reg989 = ((((reg945 ? (reg883 ^ (8'ha2)) : reg950) == ((reg980 ?
                          (8'hac) : reg956) ^~ $unsigned(wire914))) ?
                      $signed(wire869) : reg978[(4'hf):(3'h7)]) ?
                  $signed((~^((reg895 != reg948) ?
                      (!reg939) : $signed(reg902)))) : (wire869[(1'h1):(1'h0)] ?
                      $signed(reg888[(3'h5):(1'h1)]) : (reg888[(4'hc):(4'hc)] ?
                          forvar977 : $unsigned(reg917))));
            end
          else
            begin
              reg986 = (~&(|(((^wire866) || (reg956 ?
                  reg910 : reg876)) ^ (wire864[(2'h2):(1'h0)] >>> (reg986 > reg943)))));
            end
          if ({((($unsigned((7'h41)) ? $signed(reg956) : (|(8'hb0))) ?
                  reg883 : (reg873[(2'h3):(2'h3)] ?
                      (~|reg888) : (!reg918))) ^~ {reg977,
                  ($unsigned(wire912) ?
                      reg905[(1'h0):(1'h0)] : $signed((7'h46)))})})
            begin
              reg990 <= reg874[(3'h4):(3'h4)];
              reg991 <= {($signed($unsigned((wire900 ? reg910 : reg969))) ?
                      $signed($unsigned({reg962})) : reg888)};
              reg992 = $signed(($signed($unsigned((8'hb4))) <= reg887[(4'he):(4'hd)]));
            end
          else
            begin
              reg992 = (reg876[(4'ha):(4'ha)] | wire868[(4'ha):(1'h0)]);
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module709
#(parameter param820 = (^~{(|((!(7'h42)) ? ((8'h9c) ? (8'hbb) : (8'hbc)) : ((8'hab) ? (7'h41) : (7'h49)))), ((~^((8'hb6) <= (8'had))) > ((-(8'h9e)) ? ((8'hb4) ^~ (8'hb5)) : ((8'ha3) ? (8'h9d) : (8'hb2))))}))
(y, clk, wire713, wire712, wire711, wire710);
  output wire [(32'h57d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h4):(1'h0)] wire713;
  input wire [(4'hd):(1'h0)] wire712;
  input wire [(3'h6):(1'h0)] wire711;
  input wire signed [(4'h8):(1'h0)] wire710;
  reg signed [(3'h5):(1'h0)] reg819 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg817 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg816 = (1'h0);
  reg [(3'h6):(1'h0)] reg814 = (1'h0);
  reg [(2'h3):(1'h0)] reg813 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg812 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg811 = (1'h0);
  reg [(4'h9):(1'h0)] reg810 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg804 = (1'h0);
  reg [(2'h2):(1'h0)] reg803 = (1'h0);
  reg [(5'h13):(1'h0)] reg795 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg794 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg791 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg790 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg784 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg781 = (1'h0);
  reg [(5'h17):(1'h0)] reg778 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg786 = (1'h0);
  reg [(4'h9):(1'h0)] reg785 = (1'h0);
  reg [(4'he):(1'h0)] reg782 = (1'h0);
  reg [(4'h8):(1'h0)] reg779 = (1'h0);
  reg [(4'hf):(1'h0)] reg776 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg775 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg774 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg772 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg771 = (1'h0);
  reg [(5'h12):(1'h0)] reg770 = (1'h0);
  reg [(4'hf):(1'h0)] reg767 = (1'h0);
  reg [(5'h16):(1'h0)] reg763 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg760 = (1'h0);
  reg [(5'h14):(1'h0)] reg759 = (1'h0);
  reg [(4'ha):(1'h0)] reg757 = (1'h0);
  reg [(2'h3):(1'h0)] reg752 = (1'h0);
  reg [(3'h7):(1'h0)] reg751 = (1'h0);
  reg [(4'h9):(1'h0)] reg750 = (1'h0);
  reg [(5'h17):(1'h0)] reg749 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg746 = (1'h0);
  reg [(4'h9):(1'h0)] reg744 = (1'h0);
  reg [(5'h14):(1'h0)] reg743 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg742 = (1'h0);
  reg [(4'he):(1'h0)] reg739 = (1'h0);
  reg [(2'h3):(1'h0)] reg737 = (1'h0);
  reg [(5'h18):(1'h0)] reg734 = (1'h0);
  reg [(5'h18):(1'h0)] reg732 = (1'h0);
  reg [(4'h8):(1'h0)] reg731 = (1'h0);
  reg [(5'h15):(1'h0)] reg730 = (1'h0);
  reg [(4'h8):(1'h0)] reg728 = (1'h0);
  reg [(4'h8):(1'h0)] reg727 = (1'h0);
  reg [(4'hb):(1'h0)] reg725 = (1'h0);
  reg [(4'hb):(1'h0)] reg722 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg720 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg717 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg716 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg715 = (1'h0);
  reg [(4'ha):(1'h0)] reg818 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg815 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar809 = (1'h0);
  reg [(5'h10):(1'h0)] reg808 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg807 = (1'h0);
  reg [(4'he):(1'h0)] reg806 = (1'h0);
  reg [(3'h6):(1'h0)] reg805 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar802 = (1'h0);
  reg [(4'hf):(1'h0)] reg801 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg800 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar799 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg798 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar797 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg796 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg793 = (1'h0);
  reg [(5'h12):(1'h0)] reg792 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar789 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg788 = (1'h0);
  reg [(5'h12):(1'h0)] reg787 = (1'h0);
  reg [(5'h14):(1'h0)] forvar784 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg783 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar781 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg780 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar778 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg777 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg773 = (1'h0);
  reg [(4'hd):(1'h0)] reg769 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar768 = (1'h0);
  reg [(5'h17):(1'h0)] reg766 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg765 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg764 = (1'h0);
  reg [(4'he):(1'h0)] forvar762 = (1'h0);
  reg [(3'h4):(1'h0)] forvar761 = (1'h0);
  reg [(4'h9):(1'h0)] reg758 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg756 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg755 = (1'h0);
  reg [(3'h5):(1'h0)] reg754 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg753 = (1'h0);
  reg [(5'h11):(1'h0)] forvar748 = (1'h0);
  reg [(5'h17):(1'h0)] reg747 = (1'h0);
  reg [(5'h14):(1'h0)] reg748 = (1'h0);
  reg [(4'hd):(1'h0)] forvar747 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg745 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar741 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar740 = (1'h0);
  reg [(4'h8):(1'h0)] reg738 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg736 = (1'h0);
  reg [(5'h12):(1'h0)] reg735 = (1'h0);
  reg [(3'h4):(1'h0)] forvar733 = (1'h0);
  reg [(3'h7):(1'h0)] forvar729 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg726 = (1'h0);
  reg [(4'hd):(1'h0)] reg724 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar723 = (1'h0);
  reg [(4'hb):(1'h0)] reg721 = (1'h0);
  reg [(2'h2):(1'h0)] reg719 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg718 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar714 = (1'h0);
  assign y = {reg819,
                 reg817,
                 reg816,
                 reg814,
                 reg813,
                 reg812,
                 reg811,
                 reg810,
                 reg804,
                 reg803,
                 reg795,
                 reg794,
                 reg791,
                 reg790,
                 reg784,
                 reg781,
                 reg778,
                 reg786,
                 reg785,
                 reg782,
                 reg779,
                 reg776,
                 reg775,
                 reg774,
                 reg772,
                 reg771,
                 reg770,
                 reg767,
                 reg763,
                 reg760,
                 reg759,
                 reg757,
                 reg752,
                 reg751,
                 reg750,
                 reg749,
                 reg746,
                 reg744,
                 reg743,
                 reg742,
                 reg739,
                 reg737,
                 reg734,
                 reg732,
                 reg731,
                 reg730,
                 reg728,
                 reg727,
                 reg725,
                 reg722,
                 reg720,
                 reg717,
                 reg716,
                 reg715,
                 reg818,
                 reg815,
                 forvar809,
                 reg808,
                 reg807,
                 reg806,
                 reg805,
                 forvar802,
                 reg801,
                 reg800,
                 forvar799,
                 reg798,
                 forvar797,
                 reg796,
                 reg793,
                 reg792,
                 forvar789,
                 reg788,
                 reg787,
                 forvar784,
                 reg783,
                 forvar781,
                 reg780,
                 forvar778,
                 reg777,
                 reg773,
                 reg769,
                 forvar768,
                 reg766,
                 reg765,
                 reg764,
                 forvar762,
                 forvar761,
                 reg758,
                 reg756,
                 reg755,
                 reg754,
                 reg753,
                 forvar748,
                 reg747,
                 reg748,
                 forvar747,
                 reg745,
                 forvar741,
                 forvar740,
                 reg738,
                 reg736,
                 reg735,
                 forvar733,
                 forvar729,
                 reg726,
                 reg724,
                 forvar723,
                 reg721,
                 reg719,
                 reg718,
                 forvar714,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar714 = (1'h0); (forvar714 < (2'h2)); forvar714 = (forvar714 + (1'h1)))
        begin
          reg715 <= (~&({(wire710[(1'h1):(1'h1)] ^ wire710[(3'h5):(3'h5)])} >= $signed({{wire713},
              $signed((8'h9f))})));
          reg716 <= reg715[(4'h9):(2'h2)];
          if (wire710)
            begin
              reg717 <= wire712[(4'hb):(1'h0)];
              reg718 = ($unsigned((~&$signed((wire711 & wire710)))) <= (~|($signed({(8'hb5)}) ?
                  reg715[(2'h3):(1'h0)] : ((wire713 << reg715) | wire713))));
              reg719 = (wire712[(4'h8):(3'h4)] ?
                  $signed($unsigned(reg715[(4'hc):(3'h6)])) : ($signed(reg717[(1'h1):(1'h1)]) ?
                      (wire710[(2'h2):(1'h0)] ?
                          ((8'ha4) ? wire710 : (~(8'ha4))) : (wire712 ?
                              (~|reg715) : reg716[(1'h0):(1'h0)])) : reg716));
            end
          else
            begin
              reg717 <= reg717[(2'h3):(2'h2)];
            end
          reg720 <= (~&(reg716[(1'h1):(1'h1)] ?
              (~$signed(reg718[(4'ha):(4'h9)])) : ($unsigned(((7'h41) ^ reg716)) ?
                  $unsigned($unsigned(forvar714)) : (^(reg718 ?
                      (7'h49) : reg718)))));
        end
      reg721 = reg719;
      reg722 <= reg719;
    end
  always
    @(posedge clk) begin
      for (forvar723 = (1'h0); (forvar723 < (2'h3)); forvar723 = (forvar723 + (1'h1)))
        begin
          reg724 = $signed($signed(forvar723[(4'h9):(1'h0)]));
          if ($signed(($unsigned({reg715}) ?
              $signed($signed(reg724)) : (~&reg716))))
            begin
              reg725 <= ($unsigned($unsigned($unsigned(reg716))) & reg720[(3'h4):(1'h1)]);
            end
          else
            begin
              reg726 = $unsigned((~&wire710));
              reg727 <= ($unsigned(forvar723[(1'h1):(1'h0)]) ~^ (reg717 ^~ reg722));
              reg728 <= (~^($signed({reg716,
                  $unsigned(wire712)}) > wire711[(3'h6):(3'h6)]));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar729 = (1'h0); (forvar729 < (3'h4)); forvar729 = (forvar729 + (1'h1)))
        begin
          if ((-$unsigned(reg717)))
            begin
              reg730 <= (8'hb1);
            end
          else
            begin
              reg730 <= (($signed(reg722) ?
                      (^(~reg730)) : (&reg727[(2'h2):(1'h1)])) ?
                  ({$unsigned($unsigned(reg727)),
                      ({(7'h44),
                          reg727} < (~^reg727))} < {{reg716[(2'h2):(1'h1)],
                          reg722[(3'h4):(3'h4)]},
                      (^$signed(wire710))}) : $signed(reg728[(2'h2):(2'h2)]));
              reg731 <= (!wire711[(1'h1):(1'h1)]);
              reg732 <= (($unsigned((+(~|wire710))) != reg717[(2'h3):(2'h3)]) ?
                  (!{wire710}) : ({(~|reg725[(1'h1):(1'h0)])} ?
                      ({wire711, (reg720 && (8'hac))} || ((wire713 ?
                          reg727 : wire711) << reg715[(4'h9):(1'h0)])) : reg715));
            end
          for (forvar733 = (1'h0); (forvar733 < (1'h1)); forvar733 = (forvar733 + (1'h1)))
            begin
              reg734 <= ($unsigned(wire710[(4'h8):(3'h7)]) ?
                  {$unsigned($signed(reg720))} : $unsigned((reg715[(3'h7):(1'h0)] ?
                      $signed({forvar729}) : {(forvar729 || reg732)})));
              reg735 = reg725[(4'hb):(4'h8)];
              reg736 = {(&(reg716 << wire713[(1'h0):(1'h0)])),
                  ({(^reg730), reg732} ?
                      reg727 : $signed(reg727[(1'h0):(1'h0)]))};
              reg737 <= reg727;
            end
          reg738 = (-{$unsigned({$signed(reg737), reg730})});
        end
    end
  always
    @(posedge clk) begin
      reg739 <= wire710[(1'h1):(1'h0)];
      for (forvar740 = (1'h0); (forvar740 < (1'h1)); forvar740 = (forvar740 + (1'h1)))
        begin
          for (forvar741 = (1'h0); (forvar741 < (3'h4)); forvar741 = (forvar741 + (1'h1)))
            begin
              reg742 <= (reg717 + $signed($unsigned({(reg715 ?
                      forvar740 : reg725),
                  reg730})));
            end
          reg743 <= ((reg727[(1'h1):(1'h0)] ^~ $signed((reg722[(3'h4):(1'h0)] ?
                  {wire710} : (reg732 ? wire711 : reg731)))) ?
              ($unsigned($unsigned((reg737 != reg725))) >> (~&(!reg742))) : $signed(reg731[(3'h7):(3'h6)]));
          reg744 <= wire713;
        end
    end
  always
    @(posedge clk) begin
      if ($signed((+reg734)))
        begin
          reg745 = ($unsigned((reg720[(1'h0):(1'h0)] ?
              (!(reg717 ?
                  reg743 : reg725)) : $signed(reg722))) > $signed((+reg743)));
          reg746 <= (~^reg717[(2'h3):(1'h0)]);
          for (forvar747 = (1'h0); (forvar747 < (1'h0)); forvar747 = (forvar747 + (1'h1)))
            begin
              reg748 = {$unsigned({reg746, (&$signed(reg745))})};
              reg749 <= ($unsigned((((+wire711) ^ (&reg732)) <<< reg737)) ?
                  (!{reg717[(1'h0):(1'h0)],
                      wire711}) : {($signed((reg734 != (7'h45))) > {reg745,
                          reg731})});
              reg750 <= reg728[(2'h2):(2'h2)];
              reg751 <= $signed(reg743);
              reg752 <= ({$signed($signed($unsigned(wire712))),
                  wire712[(4'h9):(3'h7)]} || $unsigned({reg715, reg744}));
            end
        end
      else
        begin
          reg746 <= reg728;
          reg747 = $signed(($signed({$unsigned(reg717)}) && {(wire713[(2'h3):(1'h1)] ?
                  $signed((8'h9e)) : (reg749 <<< reg720))}));
          for (forvar748 = (1'h0); (forvar748 < (1'h0)); forvar748 = (forvar748 + (1'h1)))
            begin
              reg753 = (($unsigned(((~&forvar747) > (~reg737))) ?
                  (((^~reg730) && $signed(reg730)) ?
                      ((reg745 ? reg750 : reg715) ?
                          (reg746 && reg734) : reg737[(2'h3):(2'h2)]) : (!$unsigned(reg745))) : {forvar748[(4'ha):(1'h1)],
                      reg732}) <= (&(((reg716 ?
                      wire710 : reg727) ^ $unsigned(wire712)) ?
                  reg734 : $unsigned(wire712))));
              reg754 = $unsigned(wire711[(1'h1):(1'h1)]);
              reg755 = reg742[(3'h5):(2'h2)];
            end
          reg756 = reg742;
        end
      if (reg749[(4'hf):(4'h8)])
        begin
          reg757 <= $unsigned(reg751[(3'h5):(3'h4)]);
          reg758 = $signed(reg750[(2'h2):(1'h1)]);
        end
      else
        begin
          reg758 = reg753;
          reg759 <= reg756[(1'h0):(1'h0)];
          reg760 <= (^~$unsigned((($unsigned(reg753) ?
                  (reg737 ? reg739 : wire713) : (wire710 >= reg754)) ?
              (reg745 ?
                  (|reg757) : {reg749,
                      reg758}) : $signed(((8'ha1) < reg742)))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar761 = (1'h0); (forvar761 < (3'h4)); forvar761 = (forvar761 + (1'h1)))
        begin
          for (forvar762 = (1'h0); (forvar762 < (2'h3)); forvar762 = (forvar762 + (1'h1)))
            begin
              reg763 <= {reg727[(1'h0):(1'h0)], wire712[(4'h8):(2'h2)]};
              reg764 = reg716;
              reg765 = ($unsigned(($signed(reg742) > $unsigned(reg743[(3'h7):(3'h6)]))) >>> {$unsigned(reg757[(3'h5):(2'h3)]),
                  wire712});
            end
        end
      reg766 = (($unsigned(reg746) ?
              (($unsigned(reg751) + $unsigned(reg764)) + $unsigned($unsigned(wire712))) : (~^(8'hae))) ?
          (reg725 * reg720) : (!(reg739 ?
              ((wire712 ? reg765 : reg728) * (reg730 ?
                  reg746 : reg730)) : {{(8'haa)}})));
      reg767 <= (+reg764[(4'h9):(2'h3)]);
      for (forvar768 = (1'h0); (forvar768 < (1'h1)); forvar768 = (forvar768 + (1'h1)))
        begin
          reg769 = (|(reg763 ? $unsigned(reg751) : reg742));
          reg770 <= reg749[(3'h4):(3'h4)];
          reg771 <= $signed((|({reg717} & {(|(8'h9f)), (^~(8'ha4))})));
        end
      if ({((reg715 ?
                  (~{forvar768, reg722}) : ((reg771 & reg769) ?
                      reg731[(3'h4):(1'h1)] : (|reg725))) ?
              {$unsigned(reg731)} : $unsigned($signed(reg720)))})
        begin
          if (forvar762[(1'h0):(1'h0)])
            begin
              reg772 <= ((wire713[(1'h1):(1'h0)] == reg757) ?
                  forvar768[(1'h0):(1'h0)] : $signed((reg769 ?
                      (^(wire713 < reg725)) : forvar762)));
            end
          else
            begin
              reg773 = (8'hb5);
              reg774 <= $unsigned({(^($signed(wire713) - forvar762[(4'h9):(2'h3)]))});
              reg775 <= {reg743[(4'hd):(3'h4)]};
              reg776 <= $unsigned($unsigned($signed($signed(reg743))));
              reg777 = $unsigned(reg775);
            end
          for (forvar778 = (1'h0); (forvar778 < (1'h0)); forvar778 = (forvar778 + (1'h1)))
            begin
              reg779 <= $unsigned($signed(reg764[(4'hd):(1'h1)]));
              reg780 = $signed(reg744[(3'h4):(1'h0)]);
            end
          for (forvar781 = (1'h0); (forvar781 < (2'h2)); forvar781 = (forvar781 + (1'h1)))
            begin
              reg782 <= $unsigned(($signed($unsigned($signed(forvar762))) ?
                  $signed(reg716[(1'h0):(1'h0)]) : {forvar778[(2'h2):(2'h2)]}));
              reg783 = $signed($unsigned(((reg769[(4'h9):(3'h4)] ?
                      reg776 : reg752[(2'h2):(1'h0)]) ?
                  (~|(wire710 * reg765)) : reg771[(3'h6):(2'h2)])));
            end
          for (forvar784 = (1'h0); (forvar784 < (2'h3)); forvar784 = (forvar784 + (1'h1)))
            begin
              reg785 <= $unsigned((&($signed($signed(reg725)) - $unsigned(reg765[(3'h6):(3'h4)]))));
              reg786 <= {$signed((^{(reg752 ? reg783 : reg765)})),
                  (reg732 << $signed(((reg785 >> reg771) || (|reg772))))};
            end
        end
      else
        begin
          reg773 = reg757[(2'h2):(1'h1)];
          reg777 = $unsigned(reg780);
          if ($unsigned($unsigned($signed((reg731 ?
              $signed(reg779) : reg742)))))
            begin
              reg778 <= ({(((8'hb3) ? wire713 : $unsigned((8'hba))) ?
                          $signed((reg717 | reg751)) : ((reg760 > (7'h45)) ?
                              reg770 : (wire712 ? reg720 : reg737))),
                      (+reg779)} ?
                  reg763 : ($unsigned($signed(reg767[(3'h4):(1'h0)])) || (8'hb8)));
              reg779 <= (|((^~$signed($unsigned(reg771))) ?
                  $unsigned(({reg786, reg771} & {reg717,
                      (8'hb6)})) : (^~(&((8'hab) << wire711)))));
              reg780 = (-((reg766[(3'h5):(1'h0)] ?
                      wire710[(3'h7):(3'h7)] : (reg770[(4'hd):(2'h2)] <= reg731)) ?
                  $signed(reg778) : reg725));
              reg781 <= $signed(({{reg760}} ?
                  $signed(($signed(reg785) ?
                      $unsigned(forvar781) : $unsigned(reg732))) : reg765[(4'h9):(3'h5)]));
            end
          else
            begin
              reg778 <= reg780;
              reg779 <= reg785;
            end
          reg783 = forvar778[(3'h6):(2'h2)];
          if ($unsigned(reg766))
            begin
              reg784 <= ((-$unsigned(((~^reg732) << $signed(reg720)))) != {($unsigned($unsigned(reg725)) & forvar761),
                  reg746[(1'h1):(1'h1)]});
            end
          else
            begin
              reg784 <= reg783;
              reg787 = wire712[(3'h5):(1'h1)];
              reg788 = (((7'h46) < ((~^(reg730 ? (8'hab) : (8'ha7))) ?
                  $signed((reg722 <= reg742)) : $signed({reg764}))) <= ({((&reg744) ?
                      reg774[(4'hf):(4'h9)] : $signed(reg760)),
                  $signed(reg731)} >= $unsigned(forvar761)));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar789 = (1'h0); (forvar789 < (2'h3)); forvar789 = (forvar789 + (1'h1)))
        begin
          if (reg742[(2'h3):(2'h3)])
            begin
              reg790 <= {(wire710 ^ wire712[(2'h3):(2'h3)]),
                  ($signed(((reg728 ? wire713 : reg742) == (wire710 ?
                          reg739 : reg728))) ?
                      $signed(reg779) : reg734[(5'h12):(2'h3)])};
              reg791 <= {{((reg771 ? reg750[(4'h8):(3'h5)] : (8'h9d)) ?
                          $signed((^~reg722)) : $signed(reg737[(1'h0):(1'h0)]))}};
              reg792 = ((^~reg784[(3'h5):(1'h1)]) | {reg779[(1'h0):(1'h0)],
                  reg720[(3'h5):(1'h0)]});
              reg793 = reg722;
            end
          else
            begin
              reg792 = (-$unsigned({(reg767[(4'hd):(3'h4)] ?
                      reg772[(3'h5):(2'h2)] : $signed(reg779))}));
              reg794 <= {{{(^$unsigned(reg784))}},
                  $unsigned((&reg759[(4'h8):(4'h8)]))};
            end
          reg795 <= reg752;
          reg796 = ($unsigned(reg746[(1'h1):(1'h0)]) ^ reg715);
        end
      for (forvar797 = (1'h0); (forvar797 < (3'h4)); forvar797 = (forvar797 + (1'h1)))
        begin
          reg798 = reg770;
          for (forvar799 = (1'h0); (forvar799 < (1'h1)); forvar799 = (forvar799 + (1'h1)))
            begin
              reg800 = (|reg798[(3'h7):(3'h5)]);
              reg801 = ($unsigned(((~$signed(reg717)) ?
                      reg717 : (^~$signed(reg752)))) ?
                  ($signed((forvar789 - reg774)) << $unsigned($unsigned($signed((7'h45))))) : (^~(&reg781[(2'h2):(2'h2)])));
            end
          for (forvar802 = (1'h0); (forvar802 < (2'h2)); forvar802 = (forvar802 + (1'h1)))
            begin
              reg803 <= reg737;
              reg804 <= $signed(((reg750[(3'h5):(1'h1)] ?
                  ($unsigned(reg759) ?
                      $signed((8'ha7)) : $unsigned(reg720)) : ((reg784 << reg732) ?
                      wire712[(4'hb):(4'hb)] : $signed((7'h44)))) <= (~reg743)));
              reg805 = $signed(({({reg759} ?
                      $unsigned(reg778) : $signed(reg759)),
                  ($unsigned(reg742) >= (reg742 ?
                      reg790 : reg798))} ~^ (((~forvar799) ?
                      (reg771 ? (8'hb7) : reg795) : (~^reg795)) ?
                  (reg781 >>> reg751[(3'h5):(1'h0)]) : $unsigned((forvar789 < reg728)))));
            end
          reg806 = (reg757[(3'h7):(3'h6)] ?
              ({(~|{reg795}),
                  $unsigned($unsigned(reg785))} + reg795) : (!$signed((8'hb7))));
          reg807 = (-$signed(reg727[(3'h5):(1'h1)]));
        end
      reg808 = {$unsigned($unsigned(reg796[(1'h1):(1'h1)])), reg746};
      for (forvar809 = (1'h0); (forvar809 < (1'h1)); forvar809 = (forvar809 + (1'h1)))
        begin
          if (reg803[(1'h0):(1'h0)])
            begin
              reg810 <= (((^$unsigned($unsigned(reg795))) ?
                      $signed({(8'ha6), $signed((8'h9f))}) : {reg779,
                          ($signed(forvar802) ?
                              reg790[(2'h2):(2'h2)] : $signed(reg798))}) ?
                  (~{$unsigned(((8'ha4) ? reg763 : forvar797)),
                      reg722[(3'h4):(2'h3)]}) : wire712);
              reg811 <= ($unsigned($signed($unsigned(reg760[(2'h3):(2'h3)]))) ?
                  $unsigned(reg806[(3'h7):(1'h0)]) : $unsigned($unsigned((^~(|reg717)))));
              reg812 <= $unsigned($unsigned(reg779));
              reg813 <= $unsigned($signed((reg716[(2'h2):(1'h1)] ~^ {(8'hb3),
                  reg810[(2'h3):(1'h0)]})));
              reg814 <= $unsigned(reg734[(5'h12):(2'h2)]);
            end
          else
            begin
              reg815 = (8'ha1);
              reg816 <= $unsigned({$signed($unsigned(reg749[(4'h9):(3'h4)]))});
              reg817 <= $unsigned(((~^reg744) < (~reg790)));
              reg818 = $unsigned(($unsigned((((7'h46) ? reg794 : reg730) ?
                  $signed(reg808) : (reg759 ? reg804 : reg770))) <<< reg774));
              reg819 <= (7'h45);
            end
        end
    end
endmodule