(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h298):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire3;
  input wire [(4'hc):(1'h0)] wire2;
  input wire [(5'h11):(1'h0)] wire1;
  input wire [(5'h15):(1'h0)] wire0;
  wire [(3'h7):(1'h0)] wire641;
  wire [(3'h4):(1'h0)] wire640;
  wire signed [(2'h3):(1'h0)] wire639;
  wire [(4'he):(1'h0)] wire632;
  wire signed [(3'h4):(1'h0)] wire106;
  wire signed [(5'h15):(1'h0)] wire104;
  wire signed [(3'h7):(1'h0)] wire634;
  wire signed [(5'h11):(1'h0)] wire635;
  wire [(2'h3):(1'h0)] wire636;
  wire [(4'hb):(1'h0)] wire637;
  reg [(3'h5):(1'h0)] reg157 = (1'h0);
  reg [(4'hf):(1'h0)] reg151 = (1'h0);
  reg signed [(4'he):(1'h0)] reg149 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg148 = (1'h0);
  reg [(5'h12):(1'h0)] reg147 = (1'h0);
  reg [(4'h8):(1'h0)] reg139 = (1'h0);
  reg [(5'h10):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg131 = (1'h0);
  reg [(5'h14):(1'h0)] reg130 = (1'h0);
  reg [(5'h10):(1'h0)] reg129 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg122 = (1'h0);
  reg [(3'h6):(1'h0)] reg121 = (1'h0);
  reg [(3'h5):(1'h0)] reg118 = (1'h0);
  reg [(4'ha):(1'h0)] reg116 = (1'h0);
  reg [(4'ha):(1'h0)] reg115 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg113 = (1'h0);
  reg [(2'h3):(1'h0)] reg110 = (1'h0);
  reg [(4'ha):(1'h0)] reg108 = (1'h0);
  reg [(4'hf):(1'h0)] reg158 = (1'h0);
  reg [(5'h13):(1'h0)] reg156 = (1'h0);
  reg [(3'h7):(1'h0)] forvar155 = (1'h0);
  reg [(4'hc):(1'h0)] reg154 = (1'h0);
  reg [(2'h3):(1'h0)] forvar153 = (1'h0);
  reg [(4'hf):(1'h0)] forvar152 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg150 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg146 = (1'h0);
  reg [(5'h14):(1'h0)] reg145 = (1'h0);
  reg [(3'h6):(1'h0)] reg144 = (1'h0);
  reg [(3'h4):(1'h0)] forvar143 = (1'h0);
  reg [(5'h14):(1'h0)] reg142 = (1'h0);
  reg [(4'h9):(1'h0)] forvar141 = (1'h0);
  reg [(4'ha):(1'h0)] reg140 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg138 = (1'h0);
  reg [(4'h8):(1'h0)] forvar137 = (1'h0);
  reg [(2'h2):(1'h0)] forvar136 = (1'h0);
  reg [(2'h3):(1'h0)] reg135 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg133 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar132 = (1'h0);
  reg [(4'h8):(1'h0)] reg128 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar126 = (1'h0);
  reg [(3'h4):(1'h0)] forvar125 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg123 = (1'h0);
  reg [(4'hd):(1'h0)] reg120 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar119 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar117 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar114 = (1'h0);
  reg [(3'h5):(1'h0)] reg112 = (1'h0);
  reg [(5'h15):(1'h0)] reg111 = (1'h0);
  reg [(4'h9):(1'h0)] forvar109 = (1'h0);
  reg [(5'h14):(1'h0)] forvar107 = (1'h0);
  assign y = {wire641,
                 wire640,
                 wire639,
                 wire632,
                 wire106,
                 wire104,
                 wire634,
                 wire635,
                 wire636,
                 wire637,
                 reg157,
                 reg151,
                 reg149,
                 reg148,
                 reg147,
                 reg139,
                 reg134,
                 reg131,
                 reg130,
                 reg129,
                 reg127,
                 reg122,
                 reg121,
                 reg118,
                 reg116,
                 reg115,
                 reg113,
                 reg110,
                 reg108,
                 reg158,
                 reg156,
                 forvar155,
                 reg154,
                 forvar153,
                 forvar152,
                 reg150,
                 reg146,
                 reg145,
                 reg144,
                 forvar143,
                 reg142,
                 forvar141,
                 reg140,
                 reg138,
                 forvar137,
                 forvar136,
                 reg135,
                 reg133,
                 forvar132,
                 reg128,
                 forvar126,
                 forvar125,
                 reg124,
                 reg123,
                 reg120,
                 forvar119,
                 forvar117,
                 forvar114,
                 reg112,
                 reg111,
                 forvar109,
                 forvar107,
                 (1'h0)};
  module4 #() modinst105 (.wire6(wire2), .wire8(wire3), .wire5(wire0), .wire7(wire1), .clk(clk), .y(wire104));
  assign wire106 = $signed($signed($signed(wire2[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      for (forvar107 = (1'h0); (forvar107 < (1'h0)); forvar107 = (forvar107 + (1'h1)))
        begin
          reg108 <= $unsigned(wire2);
        end
      for (forvar109 = (1'h0); (forvar109 < (1'h1)); forvar109 = (forvar109 + (1'h1)))
        begin
          if ({$signed(((8'ha5) ? forvar107 : (~$signed(wire0))))})
            begin
              reg110 <= (wire104[(1'h1):(1'h0)] >> ((forvar107 ?
                  $unsigned({wire3, wire106}) : ((reg108 ?
                      (7'h44) : wire2) >= {reg108})) >>> (!{(~|(8'hb6))})));
              reg111 = (^~$signed($signed((&((8'hb4) ? reg110 : wire2)))));
            end
          else
            begin
              reg111 = $signed((wire104[(5'h11):(4'ha)] != ($unsigned((reg111 ?
                      wire0 : forvar107)) ?
                  reg111[(2'h2):(1'h1)] : $signed((!wire104)))));
              reg112 = wire1[(2'h2):(2'h2)];
            end
          reg113 <= {(&reg110[(2'h3):(2'h3)])};
          for (forvar114 = (1'h0); (forvar114 < (1'h0)); forvar114 = (forvar114 + (1'h1)))
            begin
              reg115 <= ($signed(wire0) <<< ((({forvar114, (8'ha0)} ?
                  forvar107[(4'hb):(1'h0)] : {reg108}) == (&reg112)) || $signed(((forvar114 ^ reg111) >> reg113))));
              reg116 <= (~{reg115, $signed($signed((!reg115)))});
            end
          for (forvar117 = (1'h0); (forvar117 < (2'h2)); forvar117 = (forvar117 + (1'h1)))
            begin
              reg118 <= ((-($signed((reg112 ?
                  wire3 : wire104)) > (-reg113[(4'hb):(4'h8)]))) <= $unsigned(($signed((wire3 ?
                      wire106 : (8'h9d))) ?
                  (~^{wire104, forvar107}) : $unsigned(reg112))));
            end
          for (forvar119 = (1'h0); (forvar119 < (1'h1)); forvar119 = (forvar119 + (1'h1)))
            begin
              reg120 = wire3;
              reg121 <= {{$unsigned(wire104[(3'h7):(3'h7)]),
                      wire104[(4'hd):(3'h5)]},
                  (~(8'hb2))};
              reg122 <= wire3;
              reg123 = (8'haa);
            end
        end
    end
  always
    @(posedge clk) begin
      reg124 = ($signed(wire106) ?
          ((~|wire104) >> $unsigned((wire0 ?
              (wire2 | wire106) : (reg116 >> (8'hbb))))) : (~|$unsigned(reg118)));
      for (forvar125 = (1'h0); (forvar125 < (2'h2)); forvar125 = (forvar125 + (1'h1)))
        begin
          for (forvar126 = (1'h0); (forvar126 < (1'h0)); forvar126 = (forvar126 + (1'h1)))
            begin
              reg127 <= $unsigned(($signed($signed($signed(reg124))) ?
                  $signed((8'hb1)) : $unsigned((^reg116[(1'h1):(1'h1)]))));
              reg128 = ((($unsigned($signed(wire104)) ?
                      reg121[(1'h0):(1'h0)] : $unsigned((forvar126 + wire3))) <<< reg124[(2'h3):(2'h2)]) ?
                  (wire2 ?
                      (8'hb9) : {$unsigned($signed(reg121))}) : ((+$unsigned($unsigned(reg113))) != wire1));
              reg129 <= (8'hbd);
              reg130 <= (wire104[(5'h11):(1'h0)] >> $signed(reg110[(2'h2):(1'h1)]));
              reg131 <= ($signed($unsigned(((reg127 ?
                  reg110 : reg127) <= $unsigned(reg118)))) == $signed(($unsigned({wire0}) ?
                  reg108[(4'ha):(1'h1)] : ($unsigned((7'h44)) + (wire3 < reg108)))));
            end
          for (forvar132 = (1'h0); (forvar132 < (1'h0)); forvar132 = (forvar132 + (1'h1)))
            begin
              reg133 = wire0;
              reg134 <= (((!{$signed(reg116),
                  forvar125[(2'h3):(1'h1)]}) ^~ ($signed((forvar125 == reg131)) ?
                  (reg118[(2'h3):(2'h3)] ?
                      (+reg116) : (reg122 ? reg128 : (8'h9f))) : ((reg133 ?
                          wire104 : wire104) ?
                      (+wire104) : $unsigned(reg116)))) == reg124);
            end
        end
      reg135 = (wire0 ~^ wire2);
      for (forvar136 = (1'h0); (forvar136 < (3'h4)); forvar136 = (forvar136 + (1'h1)))
        begin
          for (forvar137 = (1'h0); (forvar137 < (1'h1)); forvar137 = (forvar137 + (1'h1)))
            begin
              reg138 = reg134;
              reg139 <= (reg116[(3'h7):(1'h0)] != (~^(~$unsigned((reg115 ?
                  forvar137 : (8'hbe))))));
              reg140 = ((7'h43) ? $signed(reg128) : (~(7'h44)));
            end
          for (forvar141 = (1'h0); (forvar141 < (1'h0)); forvar141 = (forvar141 + (1'h1)))
            begin
              reg142 = $unsigned(forvar141[(1'h0):(1'h0)]);
            end
          for (forvar143 = (1'h0); (forvar143 < (2'h2)); forvar143 = (forvar143 + (1'h1)))
            begin
              reg144 = reg138;
              reg145 = (~^reg133[(1'h0):(1'h0)]);
              reg146 = (~^$signed((7'h44)));
              reg147 <= $unsigned(reg116[(3'h5):(2'h3)]);
              reg148 <= reg113;
            end
          if ($unsigned($signed((~&reg128))))
            begin
              reg149 <= ((&(8'ha3)) ?
                  reg121 : $signed((forvar132[(2'h2):(2'h2)] ~^ (&(^forvar125)))));
              reg150 = reg128;
            end
          else
            begin
              reg150 = ((((8'h9c) ?
                  ($signed(forvar143) ?
                      {reg150,
                          reg139} : $signed(forvar136)) : (^reg116[(3'h7):(3'h5)])) || ($signed((|(8'ha9))) ?
                  (~^(~(8'ha6))) : $signed(wire106))) == $signed((reg150 ?
                  $signed($signed(reg116)) : ({reg122, wire1} ?
                      ((7'h44) ^ forvar141) : reg138))));
              reg151 <= $signed($unsigned(reg122[(2'h3):(2'h3)]));
            end
        end
      for (forvar152 = (1'h0); (forvar152 < (2'h2)); forvar152 = (forvar152 + (1'h1)))
        begin
          for (forvar153 = (1'h0); (forvar153 < (3'h4)); forvar153 = (forvar153 + (1'h1)))
            begin
              reg154 = (forvar143 ?
                  $signed(reg135[(1'h1):(1'h1)]) : $unsigned(((reg113 ?
                          reg131[(2'h3):(1'h0)] : (reg124 ?
                              forvar126 : reg138)) ?
                      (reg142[(4'hc):(2'h2)] - $unsigned((8'ha2))) : {$signed(forvar132)})));
            end
          for (forvar155 = (1'h0); (forvar155 < (1'h1)); forvar155 = (forvar155 + (1'h1)))
            begin
              reg156 = reg108;
              reg157 <= wire1;
              reg158 = (forvar153[(2'h2):(2'h2)] ?
                  reg131[(2'h3):(2'h3)] : $unsigned((($unsigned(wire1) >> reg127[(1'h1):(1'h1)]) ?
                      {$signed(reg122),
                          (~&reg151)} : $unsigned(forvar141[(3'h5):(2'h2)]))));
            end
        end
    end
  module159 #() modinst633 (.wire163(reg149), .wire162(wire104), .wire160(reg147), .y(wire632), .clk(clk), .wire161(reg131));
  assign wire634 = (~^$unsigned(($signed((wire632 ?
                       wire632 : reg131)) <<< ((~&wire3) ?
                       {reg149, reg148} : $unsigned((8'hbe))))));
  assign wire635 = ($signed(($signed((wire104 ? reg148 : wire2)) ?
                           (~reg115) : ((~|reg118) ?
                               (8'ha1) : $unsigned(wire0)))) ?
                       (~&reg134) : reg148);
  assign wire636 = (((wire1 ?
                       reg110[(2'h3):(1'h1)] : reg134) == (~wire104)) >>> ($unsigned((reg129 ?
                       (~|reg122) : (^reg121))) && reg116));
  module374 #() modinst638 (.wire377(wire632), .wire375(wire2), .clk(clk), .wire376(reg130), .y(wire637), .wire378(wire104));
  assign wire639 = wire636[(2'h2):(1'h0)];
  assign wire640 = (~$signed((^~reg118[(3'h5):(2'h3)])));
  assign wire641 = $unsigned($signed(reg130));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module159  (y, clk, wire160, wire161, wire162, wire163);
  output wire [(32'hb3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire160;
  input wire [(5'h15):(1'h0)] wire161;
  input wire signed [(5'h15):(1'h0)] wire162;
  input wire [(4'he):(1'h0)] wire163;
  wire signed [(4'he):(1'h0)] wire630;
  wire [(5'h12):(1'h0)] wire545;
  wire signed [(5'h15):(1'h0)] wire164;
  wire signed [(5'h15):(1'h0)] wire165;
  wire signed [(5'h12):(1'h0)] wire166;
  wire [(5'h15):(1'h0)] wire290;
  wire [(5'h14):(1'h0)] wire372;
  wire [(5'h15):(1'h0)] wire460;
  wire signed [(4'hf):(1'h0)] wire462;
  wire signed [(4'h9):(1'h0)] wire543;
  assign y = {wire630,
                 wire545,
                 wire164,
                 wire165,
                 wire166,
                 wire290,
                 wire372,
                 wire460,
                 wire462,
                 wire543,
                 (1'h0)};
  assign wire164 = (wire163[(4'h8):(2'h2)] <<< $unsigned(($unsigned(wire162[(2'h3):(1'h1)]) ?
                       ($unsigned(wire160) || (wire160 * (8'hba))) : (8'haa))));
  assign wire165 = (8'hb0);
  assign wire166 = {wire160};
  module167 #() modinst291 (.wire168(wire163), .clk(clk), .wire170(wire164), .y(wire290), .wire171(wire166), .wire169(wire161));
  module292 #() modinst373 (wire372, clk, wire160, wire166, wire161, wire162);
  module374 #() modinst461 (.wire377(wire164), .wire378(wire166), .y(wire460), .wire376(wire290), .clk(clk), .wire375(wire165));
  assign wire462 = $unsigned({$unsigned({{(8'ha6), wire160},
                           {wire162, wire460}}),
                       wire460[(5'h14):(1'h0)]});
  module463 #() modinst544 (.y(wire543), .wire467(wire162), .wire465(wire160), .clk(clk), .wire466(wire372), .wire464(wire164), .wire468(wire460));
  assign wire545 = (((~^(!((8'hbb) ? wire165 : wire460))) ?
                       $unsigned(((wire161 >> (8'haa)) ?
                           $unsigned(wire165) : wire460)) : wire165) || ($unsigned($unsigned($signed(wire164))) ?
                       {(8'hb6)} : $unsigned(($signed(wire165) ?
                           (&wire164) : wire163))));
  module546 #() modinst631 (wire630, clk, wire161, wire543, wire290, wire460);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module4
#(parameter param102 = (&(((&((8'hb9) ? (8'ha1) : (8'ha1))) ? (8'h9f) : (~|(|(8'had)))) ? (|(((8'ha2) ? (8'hb3) : (8'ha1)) ? {(7'h40)} : (~&(8'h9c)))) : ((~&(|(8'haf))) ? (^~((8'ha8) <<< (7'h43))) : ((~|(7'h41)) <<< (!(8'haf)))))), 
parameter param103 = (^(({((8'ha6) >= param102)} + {{param102}, ((8'h9f) ? param102 : param102)}) * {param102})))
(y, clk, wire8, wire7, wire6, wire5);
  output wire [(32'heb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hc):(1'h0)] wire8;
  input wire signed [(5'h11):(1'h0)] wire7;
  input wire [(3'h7):(1'h0)] wire6;
  input wire signed [(5'h15):(1'h0)] wire5;
  wire [(5'h11):(1'h0)] wire101;
  wire signed [(3'h6):(1'h0)] wire99;
  wire [(4'ha):(1'h0)] wire10;
  wire signed [(4'h8):(1'h0)] wire9;
  reg [(5'h13):(1'h0)] reg13 = (1'h0);
  reg [(4'ha):(1'h0)] reg14 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg16 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg17 = (1'h0);
  reg [(5'h11):(1'h0)] reg19 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg20 = (1'h0);
  reg [(5'h10):(1'h0)] reg22 = (1'h0);
  reg [(4'hb):(1'h0)] reg23 = (1'h0);
  reg [(5'h14):(1'h0)] reg25 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg26 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar24 = (1'h0);
  reg [(3'h5):(1'h0)] reg21 = (1'h0);
  reg [(5'h14):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar15 = (1'h0);
  reg [(2'h3):(1'h0)] forvar12 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar11 = (1'h0);
  assign y = {wire101,
                 wire99,
                 wire10,
                 wire9,
                 reg13,
                 reg14,
                 reg16,
                 reg17,
                 reg19,
                 reg20,
                 reg22,
                 reg23,
                 reg25,
                 reg26,
                 forvar24,
                 reg21,
                 reg18,
                 forvar15,
                 forvar12,
                 forvar11,
                 (1'h0)};
  assign wire9 = $signed(($signed(((+wire6) ?
                         $signed(wire6) : wire7[(3'h7):(3'h7)])) ?
                     (wire8 ?
                         ($signed(wire6) ?
                             {wire5} : (wire5 ?
                                 wire7 : wire5)) : ((&wire6) <<< ((8'hb9) ?
                             wire8 : wire6))) : wire5[(2'h2):(2'h2)]));
  assign wire10 = $unsigned((!$signed(wire5)));
  always
    @(posedge clk) begin
      for (forvar11 = (1'h0); (forvar11 < (2'h3)); forvar11 = (forvar11 + (1'h1)))
        begin
          for (forvar12 = (1'h0); (forvar12 < (3'h4)); forvar12 = (forvar12 + (1'h1)))
            begin
              reg13 <= wire6;
              reg14 <= $unsigned((~&{{(wire8 ? (8'ha3) : reg13)}}));
            end
          for (forvar15 = (1'h0); (forvar15 < (1'h0)); forvar15 = (forvar15 + (1'h1)))
            begin
              reg16 <= ((~|wire9) ?
                  $unsigned((^{(+wire5),
                      wire9})) : $unsigned(forvar15[(5'h11):(3'h6)]));
              reg17 <= wire7[(4'hf):(4'hc)];
              reg18 = $unsigned(wire8);
              reg19 <= reg18[(4'h8):(3'h4)];
              reg20 <= $signed(forvar11);
            end
          reg21 = $signed((~|$signed((~$unsigned(forvar15)))));
        end
      reg22 <= (wire5 ?
          ((reg21 + forvar12) ?
              $unsigned({reg14[(3'h6):(3'h6)]}) : reg18) : ((reg14 <= wire6) & $signed($unsigned(wire10))));
      reg23 <= ($signed(({((8'hb9) ? wire9 : reg19),
          wire9} <= $unsigned((8'hb6)))) ~^ (reg17[(3'h4):(1'h0)] >= (reg16[(2'h3):(2'h2)] ?
          {(reg14 ^~ wire8), $unsigned(reg16)} : $unsigned(((7'h44) ?
              (8'hbe) : (8'hba))))));
      for (forvar24 = (1'h0); (forvar24 < (3'h4)); forvar24 = (forvar24 + (1'h1)))
        begin
          reg25 <= $signed(forvar12);
        end
      reg26 = reg25[(1'h0):(1'h0)];
    end
  module27 #() modinst100 (.wire30(reg22), .clk(clk), .wire29(wire10), .y(wire99), .wire31(reg17), .wire32(wire8), .wire28(reg25));
  assign wire101 = wire10;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module27
#(parameter param97 = ((^~(+(8'hb3))) || (~^{(8'hbf), (((8'hb6) == (8'hbd)) || ((8'h9f) ? (8'hb8) : (7'h41)))})), 
parameter param98 = (!{param97, {param97}}))
(y, clk, wire32, wire31, wire30, wire29, wire28);
  output wire [(32'h2ec):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hc):(1'h0)] wire32;
  input wire [(4'hc):(1'h0)] wire31;
  input wire [(2'h2):(1'h0)] wire30;
  input wire signed [(4'h9):(1'h0)] wire29;
  input wire [(5'h14):(1'h0)] wire28;
  wire signed [(4'hd):(1'h0)] wire96;
  wire signed [(3'h5):(1'h0)] wire95;
  wire signed [(4'hb):(1'h0)] wire94;
  wire signed [(3'h5):(1'h0)] wire93;
  wire signed [(5'h13):(1'h0)] wire62;
  wire [(2'h3):(1'h0)] wire61;
  wire signed [(4'hf):(1'h0)] wire60;
  wire [(4'h8):(1'h0)] wire59;
  wire signed [(4'h9):(1'h0)] wire58;
  wire [(5'h10):(1'h0)] wire57;
  wire signed [(3'h5):(1'h0)] wire56;
  wire [(4'hc):(1'h0)] wire55;
  wire signed [(2'h2):(1'h0)] wire54;
  wire [(4'hb):(1'h0)] wire53;
  wire [(5'h13):(1'h0)] wire52;
  wire signed [(5'h10):(1'h0)] wire51;
  wire signed [(4'hc):(1'h0)] wire50;
  wire signed [(4'ha):(1'h0)] wire36;
  wire [(5'h12):(1'h0)] wire35;
  wire signed [(4'he):(1'h0)] wire34;
  wire [(3'h6):(1'h0)] wire33;
  reg [(4'h9):(1'h0)] reg92 = (1'h0);
  reg [(4'hb):(1'h0)] reg87 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg86 = (1'h0);
  reg [(4'hc):(1'h0)] reg84 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg82 = (1'h0);
  reg [(5'h14):(1'h0)] reg77 = (1'h0);
  reg [(3'h6):(1'h0)] reg75 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg73 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg71 = (1'h0);
  reg [(4'hf):(1'h0)] reg69 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg64 = (1'h0);
  reg [(4'ha):(1'h0)] reg45 = (1'h0);
  reg [(4'hd):(1'h0)] reg38 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg49 = (1'h0);
  reg [(2'h2):(1'h0)] reg48 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg47 = (1'h0);
  reg [(4'h8):(1'h0)] reg46 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg44 = (1'h0);
  reg [(3'h4):(1'h0)] reg41 = (1'h0);
  reg [(3'h7):(1'h0)] reg39 = (1'h0);
  reg [(4'hf):(1'h0)] reg37 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg91 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar90 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg89 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg88 = (1'h0);
  reg [(3'h6):(1'h0)] forvar85 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg83 = (1'h0);
  reg [(4'hb):(1'h0)] reg81 = (1'h0);
  reg [(4'hb):(1'h0)] reg80 = (1'h0);
  reg [(5'h12):(1'h0)] reg79 = (1'h0);
  reg [(2'h3):(1'h0)] forvar78 = (1'h0);
  reg signed [(4'he):(1'h0)] reg76 = (1'h0);
  reg [(2'h2):(1'h0)] forvar74 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar72 = (1'h0);
  reg [(4'h9):(1'h0)] reg70 = (1'h0);
  reg [(4'h9):(1'h0)] reg68 = (1'h0);
  reg [(2'h3):(1'h0)] forvar67 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg66 = (1'h0);
  reg [(4'hb):(1'h0)] forvar65 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar63 = (1'h0);
  reg [(2'h2):(1'h0)] reg42 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar40 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar37 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar45 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg43 = (1'h0);
  reg [(5'h13):(1'h0)] forvar42 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg40 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar38 = (1'h0);
  assign y = {wire96,
                 wire95,
                 wire94,
                 wire93,
                 wire62,
                 wire61,
                 wire60,
                 wire59,
                 wire58,
                 wire57,
                 wire56,
                 wire55,
                 wire54,
                 wire53,
                 wire52,
                 wire51,
                 wire50,
                 wire36,
                 wire35,
                 wire34,
                 wire33,
                 reg92,
                 reg87,
                 reg86,
                 reg84,
                 reg82,
                 reg77,
                 reg75,
                 reg73,
                 reg71,
                 reg69,
                 reg64,
                 reg45,
                 reg38,
                 reg49,
                 reg48,
                 reg47,
                 reg46,
                 reg44,
                 reg41,
                 reg39,
                 reg37,
                 reg91,
                 forvar90,
                 reg89,
                 reg88,
                 forvar85,
                 reg83,
                 reg81,
                 reg80,
                 reg79,
                 forvar78,
                 reg76,
                 forvar74,
                 forvar72,
                 reg70,
                 reg68,
                 forvar67,
                 reg66,
                 forvar65,
                 forvar63,
                 reg42,
                 forvar40,
                 forvar37,
                 forvar45,
                 reg43,
                 forvar42,
                 reg40,
                 forvar38,
                 (1'h0)};
  assign wire33 = (($unsigned((wire30[(1'h1):(1'h0)] ?
                          $unsigned((8'hb6)) : $signed(wire31))) ?
                      (^(((7'h40) && wire32) ^~ (~&wire29))) : (+wire31[(3'h4):(2'h3)])) >>> $signed((8'ha5)));
  assign wire34 = {(~&$unsigned(($unsigned(wire32) >> (wire32 * wire32)))),
                      (wire30 ? wire32[(4'hb):(3'h7)] : (8'hb5))};
  assign wire35 = (wire29[(3'h6):(2'h2)] ? wire28 : wire29[(3'h5):(2'h3)]);
  assign wire36 = ((wire32 - (((wire33 == wire30) ?
                          wire35 : (wire34 ~^ wire33)) ?
                      $unsigned((^wire31)) : (+((8'hb7) & wire33)))) <= {wire32,
                      (~&wire30)});
  always
    @(posedge clk) begin
      if (wire28[(4'he):(2'h2)])
        begin
          reg37 <= wire31[(2'h3):(1'h0)];
          for (forvar38 = (1'h0); (forvar38 < (2'h2)); forvar38 = (forvar38 + (1'h1)))
            begin
              reg39 <= ({(|{(^~wire28)})} ?
                  $unsigned($signed((~|wire29))) : (({(wire29 + wire30)} + $signed((!wire34))) ?
                      wire29[(3'h5):(3'h4)] : (^wire35)));
              reg40 = (+wire31[(1'h0):(1'h0)]);
              reg41 <= $unsigned($unsigned((8'hb3)));
            end
          for (forvar42 = (1'h0); (forvar42 < (1'h0)); forvar42 = (forvar42 + (1'h1)))
            begin
              reg43 = $unsigned((|($unsigned((8'hbf)) ?
                  (|(~reg37)) : {(reg40 ? wire31 : reg40)})));
              reg44 <= $signed($signed((^~(8'ha1))));
            end
          for (forvar45 = (1'h0); (forvar45 < (2'h3)); forvar45 = (forvar45 + (1'h1)))
            begin
              reg46 <= ($unsigned(reg39) ^~ (8'hbc));
              reg47 <= reg39;
              reg48 <= (8'ha5);
              reg49 <= {(wire29 ?
                      $unsigned($unsigned($signed(forvar45))) : reg48[(2'h2):(1'h1)]),
                  wire30[(1'h1):(1'h0)]};
            end
        end
      else
        begin
          for (forvar37 = (1'h0); (forvar37 < (1'h1)); forvar37 = (forvar37 + (1'h1)))
            begin
              reg38 <= (+(+(({(8'hae), reg47} ?
                  ((8'hb9) - wire35) : (wire33 ^~ (8'ha9))) ~^ $unsigned({wire33}))));
              reg39 <= wire31;
            end
          for (forvar40 = (1'h0); (forvar40 < (3'h4)); forvar40 = (forvar40 + (1'h1)))
            begin
              reg42 = {(-((~&reg49[(5'h14):(5'h10)]) ?
                      {$unsigned(reg47)} : ($unsigned(reg43) - wire33[(1'h0):(1'h0)]))),
                  $signed($unsigned((~$unsigned(reg38))))};
              reg43 = $signed(reg41);
              reg44 <= (reg46[(3'h7):(1'h0)] ^ (($unsigned((reg47 > wire31)) != wire30[(2'h2):(2'h2)]) >= forvar40[(4'h8):(1'h1)]));
              reg45 <= $signed((!$signed(wire35)));
              reg46 <= {((((^forvar37) <<< (forvar37 ? reg37 : forvar45)) ?
                      $signed($signed(wire36)) : ((+reg48) >>> (~&(8'hbb)))) && (~&((-wire34) ?
                      $signed(reg38) : {reg43, forvar45})))};
            end
        end
    end
  assign wire50 = $unsigned(($signed(((^wire28) >= (reg41 ? (7'h44) : reg46))) ?
                      reg39 : (^(+((8'ha1) * (8'had))))));
  assign wire51 = (|{(^{(reg48 ? wire30 : (8'hb9)), reg45[(1'h1):(1'h0)]}),
                      reg37});
  assign wire52 = {(+reg49[(4'hc):(3'h6)]), wire28[(3'h7):(3'h7)]};
  assign wire53 = (~(~((wire30 > (wire52 ?
                      reg48 : reg41)) & ((wire33 + (7'h44)) ?
                      reg41 : {wire34}))));
  assign wire54 = {($unsigned((~^{wire33})) * {reg46[(3'h5):(2'h2)]}),
                      $unsigned($unsigned(reg45))};
  assign wire55 = $signed(reg41);
  assign wire56 = wire32[(2'h3):(2'h2)];
  assign wire57 = ((|(($signed(wire50) ?
                          $unsigned(reg48) : (reg48 ? wire36 : wire31)) ?
                      (reg45 ?
                          reg49[(4'h9):(3'h5)] : wire50[(4'ha):(3'h5)]) : ((wire54 | wire50) - (~reg46)))) + $signed((({wire35,
                          wire31} ?
                      (reg37 < (8'hac)) : (+(8'hb6))) < (7'h44))));
  assign wire58 = ((8'hac) && $signed($unsigned(wire32[(4'h9):(4'h8)])));
  assign wire59 = ({(~&(8'h9f)), ($unsigned(wire50) + (|(+wire56)))} ?
                      (~reg37) : {reg39[(2'h2):(1'h0)]});
  assign wire60 = (reg44[(2'h2):(1'h0)] ?
                      $unsigned((^~wire55)) : wire56[(3'h4):(2'h3)]);
  assign wire61 = wire36;
  assign wire62 = (!(~^({(reg38 <<< wire57)} >> ((reg46 | wire35) ?
                      (reg38 >= (8'hbc)) : (+reg47)))));
  always
    @(posedge clk) begin
      for (forvar63 = (1'h0); (forvar63 < (2'h3)); forvar63 = (forvar63 + (1'h1)))
        begin
          reg64 <= {(reg46[(3'h4):(1'h0)] ?
                  wire36[(4'h8):(2'h2)] : (-{$signed(wire32),
                      (reg38 ? wire36 : reg46)})),
              ($unsigned(($unsigned((8'hac)) >= (~^reg37))) ?
                  (8'hbd) : ((^~(wire31 - reg49)) < ($unsigned((7'h44)) > {wire55,
                      reg49})))};
          for (forvar65 = (1'h0); (forvar65 < (1'h1)); forvar65 = (forvar65 + (1'h1)))
            begin
              reg66 = $signed((($signed(wire55) ?
                      forvar63[(4'h8):(3'h4)] : {$signed(wire54),
                          (wire31 ? wire33 : reg41)}) ?
                  (!(7'h42)) : ($signed((wire59 ?
                      wire55 : wire54)) != (~(wire36 ? wire58 : wire60)))));
            end
          for (forvar67 = (1'h0); (forvar67 < (1'h0)); forvar67 = (forvar67 + (1'h1)))
            begin
              reg68 = (^~(~^wire30[(1'h0):(1'h0)]));
              reg69 <= wire54[(1'h1):(1'h0)];
              reg70 = reg68[(1'h0):(1'h0)];
            end
          reg71 <= reg70;
        end
      for (forvar72 = (1'h0); (forvar72 < (2'h3)); forvar72 = (forvar72 + (1'h1)))
        begin
          reg73 <= (^~($unsigned((!{wire36})) ?
              (((^reg69) ? (wire58 - wire53) : {reg66, forvar63}) ?
                  (wire32 ?
                      (wire32 ?
                          wire53 : wire59) : (wire61 < wire56)) : (~^(^~forvar67))) : $signed(wire57[(3'h4):(2'h3)])));
          for (forvar74 = (1'h0); (forvar74 < (1'h0)); forvar74 = (forvar74 + (1'h1)))
            begin
              reg75 <= $unsigned($unsigned(((8'hab) - (((8'hb1) ?
                  (7'h41) : reg45) | forvar72[(4'hb):(4'h9)]))));
              reg76 = $signed({(((forvar67 ?
                      reg73 : wire62) + $signed((8'ha1))) <= wire28[(4'ha):(3'h5)])});
            end
          reg77 <= reg37;
          for (forvar78 = (1'h0); (forvar78 < (3'h4)); forvar78 = (forvar78 + (1'h1)))
            begin
              reg79 = (wire52[(3'h6):(3'h4)] + wire55);
              reg80 = wire32[(3'h4):(1'h0)];
              reg81 = ((&(~|wire36)) ? wire34[(4'hb):(4'h9)] : wire33);
              reg82 <= {reg47[(3'h4):(1'h0)]};
              reg83 = $unsigned($signed((~|(((8'hb7) && reg68) == wire30[(1'h1):(1'h1)]))));
            end
          reg84 <= forvar74;
        end
      if ((~^(!reg41)))
        begin
          for (forvar85 = (1'h0); (forvar85 < (1'h1)); forvar85 = (forvar85 + (1'h1)))
            begin
              reg86 <= wire56;
            end
          reg87 <= $signed((8'h9d));
        end
      else
        begin
          for (forvar85 = (1'h0); (forvar85 < (2'h2)); forvar85 = (forvar85 + (1'h1)))
            begin
              reg86 <= wire31[(2'h3):(2'h3)];
              reg88 = $unsigned((8'hab));
            end
          reg89 = $unsigned((reg83[(5'h10):(3'h4)] ~^ reg69));
          for (forvar90 = (1'h0); (forvar90 < (2'h3)); forvar90 = (forvar90 + (1'h1)))
            begin
              reg91 = (+reg79[(4'hc):(3'h5)]);
              reg92 <= {(+((8'hae) ? forvar67[(1'h0):(1'h0)] : reg82)),
                  ((~$signed(reg82)) ?
                      wire35[(3'h7):(3'h5)] : (+$signed($signed(forvar63))))};
            end
        end
    end
  assign wire93 = $signed((8'hb1));
  assign wire94 = $signed((!wire58[(3'h6):(1'h0)]));
  assign wire95 = $unsigned(wire55);
  assign wire96 = $unsigned((-({(reg82 | wire28), (!reg87)} ?
                      (+reg71[(5'h11):(4'hb)]) : ($unsigned((8'ha3)) > $unsigned(wire34)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module546  (y, clk, wire550, wire549, wire548, wire547);
  output wire [(32'h3aa):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h13):(1'h0)] wire550;
  input wire signed [(2'h3):(1'h0)] wire549;
  input wire signed [(4'h8):(1'h0)] wire548;
  input wire [(4'hb):(1'h0)] wire547;
  wire signed [(5'h13):(1'h0)] wire629;
  wire [(3'h7):(1'h0)] wire628;
  wire [(5'h13):(1'h0)] wire627;
  wire signed [(3'h5):(1'h0)] wire626;
  wire signed [(4'h8):(1'h0)] wire583;
  wire [(4'h9):(1'h0)] wire582;
  wire [(4'he):(1'h0)] wire571;
  wire [(5'h10):(1'h0)] wire570;
  wire [(5'h14):(1'h0)] wire569;
  wire signed [(4'h9):(1'h0)] wire568;
  wire [(3'h5):(1'h0)] wire567;
  wire signed [(5'h12):(1'h0)] wire566;
  wire [(4'hc):(1'h0)] wire555;
  wire [(4'hd):(1'h0)] wire554;
  wire signed [(4'hb):(1'h0)] wire553;
  wire [(3'h6):(1'h0)] wire552;
  wire signed [(4'hc):(1'h0)] wire551;
  reg signed [(5'h15):(1'h0)] reg625 = (1'h0);
  reg [(2'h3):(1'h0)] reg623 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg618 = (1'h0);
  reg [(4'he):(1'h0)] reg614 = (1'h0);
  reg [(3'h6):(1'h0)] reg612 = (1'h0);
  reg [(3'h5):(1'h0)] reg608 = (1'h0);
  reg [(3'h6):(1'h0)] reg607 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg606 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg604 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg601 = (1'h0);
  reg [(4'he):(1'h0)] reg599 = (1'h0);
  reg [(5'h13):(1'h0)] reg598 = (1'h0);
  reg [(5'h13):(1'h0)] reg595 = (1'h0);
  reg [(4'hf):(1'h0)] reg594 = (1'h0);
  reg [(4'he):(1'h0)] reg592 = (1'h0);
  reg [(4'hf):(1'h0)] reg589 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg588 = (1'h0);
  reg [(5'h13):(1'h0)] reg581 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg580 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg577 = (1'h0);
  reg [(5'h14):(1'h0)] reg565 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg562 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg561 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg558 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar622 = (1'h0);
  reg [(2'h2):(1'h0)] forvar621 = (1'h0);
  reg [(5'h12):(1'h0)] reg620 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg619 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg617 = (1'h0);
  reg [(4'hf):(1'h0)] reg616 = (1'h0);
  reg [(2'h3):(1'h0)] reg615 = (1'h0);
  reg [(2'h2):(1'h0)] reg613 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg611 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg610 = (1'h0);
  reg [(5'h14):(1'h0)] forvar609 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg605 = (1'h0);
  reg [(4'ha):(1'h0)] forvar603 = (1'h0);
  reg [(3'h7):(1'h0)] reg602 = (1'h0);
  reg [(2'h2):(1'h0)] reg600 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar597 = (1'h0);
  reg [(4'hd):(1'h0)] reg596 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg593 = (1'h0);
  reg [(3'h7):(1'h0)] forvar591 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar590 = (1'h0);
  reg [(3'h7):(1'h0)] reg587 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar586 = (1'h0);
  reg [(4'h9):(1'h0)] forvar585 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg584 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar579 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg578 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar576 = (1'h0);
  reg [(4'he):(1'h0)] reg575 = (1'h0);
  reg [(4'hd):(1'h0)] forvar574 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar573 = (1'h0);
  reg [(5'h12):(1'h0)] reg572 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg564 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar563 = (1'h0);
  reg [(4'h9):(1'h0)] reg560 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg559 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar557 = (1'h0);
  reg [(2'h3):(1'h0)] forvar556 = (1'h0);
  assign y = {wire629,
                 wire628,
                 wire627,
                 wire626,
                 wire583,
                 wire582,
                 wire571,
                 wire570,
                 wire569,
                 wire568,
                 wire567,
                 wire566,
                 wire555,
                 wire554,
                 wire553,
                 wire552,
                 wire551,
                 reg625,
                 reg623,
                 reg618,
                 reg614,
                 reg612,
                 reg608,
                 reg607,
                 reg606,
                 reg604,
                 reg601,
                 reg599,
                 reg598,
                 reg595,
                 reg594,
                 reg592,
                 reg589,
                 reg588,
                 reg581,
                 reg580,
                 reg577,
                 reg565,
                 reg562,
                 reg561,
                 reg558,
                 reg624,
                 forvar622,
                 forvar621,
                 reg620,
                 reg619,
                 reg617,
                 reg616,
                 reg615,
                 reg613,
                 reg611,
                 reg610,
                 forvar609,
                 reg605,
                 forvar603,
                 reg602,
                 reg600,
                 forvar597,
                 reg596,
                 reg593,
                 forvar591,
                 forvar590,
                 reg587,
                 forvar586,
                 forvar585,
                 reg584,
                 forvar579,
                 reg578,
                 forvar576,
                 reg575,
                 forvar574,
                 forvar573,
                 reg572,
                 reg564,
                 forvar563,
                 reg560,
                 reg559,
                 forvar557,
                 forvar556,
                 (1'h0)};
  assign wire551 = $signed(wire549[(1'h0):(1'h0)]);
  assign wire552 = wire551;
  assign wire553 = wire551;
  assign wire554 = wire551[(1'h0):(1'h0)];
  assign wire555 = wire551;
  always
    @(posedge clk) begin
      for (forvar556 = (1'h0); (forvar556 < (1'h1)); forvar556 = (forvar556 + (1'h1)))
        begin
          for (forvar557 = (1'h0); (forvar557 < (1'h1)); forvar557 = (forvar557 + (1'h1)))
            begin
              reg558 <= (((8'ha2) ? (+wire548) : wire551[(4'h9):(3'h7)]) ?
                  (8'hbf) : $unsigned((+wire548)));
              reg559 = wire551[(3'h6):(2'h3)];
              reg560 = ($unsigned((wire547[(2'h2):(1'h1)] >> ({wire550} >> (wire553 ?
                      (8'hb6) : forvar556)))) ?
                  (($signed(wire553) ?
                          wire550[(1'h0):(1'h0)] : $unsigned({(8'hab),
                              wire547})) ?
                      $unsigned((^$unsigned(forvar556))) : $unsigned(((8'h9c) ?
                          (wire548 <<< forvar557) : (~^(8'had))))) : $unsigned((8'h9c)));
              reg561 <= wire551[(3'h5):(1'h1)];
            end
          reg562 <= wire552[(2'h3):(1'h0)];
          for (forvar563 = (1'h0); (forvar563 < (2'h3)); forvar563 = (forvar563 + (1'h1)))
            begin
              reg564 = $unsigned(reg562);
              reg565 <= (&($unsigned(reg560) ?
                  (~^$signed((8'ha7))) : reg560[(3'h7):(3'h6)]));
            end
        end
    end
  assign wire566 = ($unsigned($signed(((&wire554) + {(8'ha0)}))) || wire547[(4'h8):(3'h6)]);
  assign wire567 = wire566[(4'h9):(1'h0)];
  assign wire568 = (^{reg562[(2'h2):(1'h1)]});
  assign wire569 = ((~wire551[(1'h1):(1'h0)]) ?
                       $signed(reg562[(3'h4):(2'h2)]) : (-((!wire547) ?
                           ((wire551 ? reg561 : (8'haf)) ?
                               {reg558,
                                   (8'hb5)} : (wire548 != wire550)) : (wire551[(4'ha):(4'ha)] ?
                               $unsigned((8'hbb)) : (wire566 <<< reg565)))));
  assign wire570 = $signed((({$unsigned(reg562),
                           reg558[(3'h7):(2'h3)]} * wire547[(3'h4):(1'h1)]) ?
                       ((wire569 ? {wire552, wire568} : $signed(wire549)) ?
                           wire548 : {(8'hbd)}) : $unsigned((wire552[(3'h4):(2'h3)] <= wire567))));
  assign wire571 = (!wire547);
  always
    @(posedge clk) begin
      reg572 = ($unsigned((8'hba)) ~^ $unsigned($unsigned(wire570[(4'hb):(3'h5)])));
    end
  always
    @(posedge clk) begin
      for (forvar573 = (1'h0); (forvar573 < (3'h4)); forvar573 = (forvar573 + (1'h1)))
        begin
          for (forvar574 = (1'h0); (forvar574 < (2'h2)); forvar574 = (forvar574 + (1'h1)))
            begin
              reg575 = $signed(((8'ha3) ^ reg558[(3'h6):(1'h1)]));
            end
          for (forvar576 = (1'h0); (forvar576 < (3'h4)); forvar576 = (forvar576 + (1'h1)))
            begin
              reg577 <= ((($unsigned(((8'hbe) ?
                      forvar573 : reg575)) <= (~(wire550 ?
                      wire550 : (8'ha5)))) ?
                  ((|(reg561 > reg561)) ?
                      ($signed(wire554) ?
                          $signed(reg561) : wire566) : (forvar573[(1'h0):(1'h0)] == wire571[(1'h0):(1'h0)])) : (forvar574 ^~ wire567[(2'h3):(2'h3)])) <<< $unsigned({wire571[(2'h3):(2'h2)],
                  (&(reg561 ? (8'ha8) : wire571))}));
            end
          reg578 = ($unsigned({$signed(wire568)}) ?
              (+$signed((+wire568))) : (reg561 + (^~(~&(reg562 ~^ (8'hbe))))));
          for (forvar579 = (1'h0); (forvar579 < (2'h3)); forvar579 = (forvar579 + (1'h1)))
            begin
              reg580 <= $signed({reg558});
              reg581 <= wire568;
            end
        end
    end
  assign wire582 = wire568[(3'h7):(3'h5)];
  assign wire583 = wire553[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg584 = $signed({wire570,
          $signed((wire551[(4'hc):(1'h1)] ?
              (wire566 >= wire566) : (wire548 != wire552)))});
      for (forvar585 = (1'h0); (forvar585 < (3'h4)); forvar585 = (forvar585 + (1'h1)))
        begin
          for (forvar586 = (1'h0); (forvar586 < (2'h2)); forvar586 = (forvar586 + (1'h1)))
            begin
              reg587 = {(reg561[(2'h3):(1'h0)] ?
                      wire571[(3'h7):(3'h4)] : {(~|(wire568 ?
                              (8'hb4) : (8'h9c))),
                          wire549[(2'h2):(1'h1)]})};
              reg588 <= (($signed($signed((&wire547))) > wire554) ^~ ((wire551 ?
                      (|wire554[(4'hb):(4'hb)]) : $signed($signed(reg584))) ?
                  (((reg558 && wire568) * $signed(wire571)) <= {reg587}) : $signed($signed(forvar585[(2'h3):(1'h0)]))));
              reg589 <= wire549;
            end
        end
      for (forvar590 = (1'h0); (forvar590 < (1'h0)); forvar590 = (forvar590 + (1'h1)))
        begin
          for (forvar591 = (1'h0); (forvar591 < (2'h2)); forvar591 = (forvar591 + (1'h1)))
            begin
              reg592 <= $signed(reg580);
              reg593 = $signed($signed(wire571[(4'he):(3'h5)]));
              reg594 <= wire569[(2'h2):(1'h1)];
              reg595 <= (8'h9f);
              reg596 = (-wire568[(1'h1):(1'h0)]);
            end
        end
      for (forvar597 = (1'h0); (forvar597 < (2'h2)); forvar597 = (forvar597 + (1'h1)))
        begin
          if ((~$unsigned((((wire566 ? reg594 : (8'h9e)) ?
              wire552 : wire552) << ((~^reg589) - $unsigned(wire571))))))
            begin
              reg598 <= ($signed((^~$unsigned((reg593 ?
                  wire566 : wire555)))) && (~^$signed($signed(reg577))));
              reg599 <= reg565[(5'h11):(4'hd)];
              reg600 = $signed($unsigned(((~|$signed((8'ha5))) ?
                  $signed((forvar585 ?
                      reg565 : reg596)) : $unsigned((^forvar591)))));
              reg601 <= (~&wire548[(3'h7):(1'h1)]);
            end
          else
            begin
              reg598 <= reg588[(3'h7):(2'h3)];
              reg600 = reg601;
              reg601 <= {$signed(reg595[(5'h11):(1'h1)]),
                  $unsigned($unsigned((-(reg581 == wire548))))};
              reg602 = (~forvar585[(2'h2):(1'h0)]);
            end
          for (forvar603 = (1'h0); (forvar603 < (1'h0)); forvar603 = (forvar603 + (1'h1)))
            begin
              reg604 <= ($signed(reg562) ?
                  (+(reg580[(3'h5):(3'h4)] << (~^$unsigned(reg562)))) : $signed((~^({wire569,
                          forvar585} ?
                      $signed(reg562) : {forvar590, reg594}))));
              reg605 = (^~wire553);
              reg606 <= {{reg589, wire551[(3'h4):(1'h1)]},
                  $unsigned((($signed(reg561) == {reg561,
                      forvar585}) | forvar585[(2'h3):(2'h3)]))};
              reg607 <= $unsigned(reg606);
            end
          reg608 <= (8'hbf);
          for (forvar609 = (1'h0); (forvar609 < (1'h1)); forvar609 = (forvar609 + (1'h1)))
            begin
              reg610 = (~|(wire553 ?
                  {(7'h41), (!(wire549 ? reg581 : wire547))} : ((8'haa) ?
                      $signed($unsigned(reg587)) : $signed($unsigned(forvar590)))));
              reg611 = $unsigned(({{(~reg587), forvar585[(4'h9):(1'h0)]},
                      ({wire570, reg588} ?
                          (reg608 ? wire566 : reg588) : $unsigned(reg584))} ?
                  (((+wire550) ^~ (-(8'hbe))) >= (~&$unsigned(forvar597))) : $unsigned(((reg558 >>> reg589) + reg604[(1'h0):(1'h0)]))));
              reg612 <= $unsigned(wire583[(1'h1):(1'h0)]);
              reg613 = ($signed((~&($unsigned(reg561) * $signed((8'hb8))))) ?
                  $unsigned((($unsigned((8'hb3)) >>> wire552[(1'h1):(1'h1)]) ?
                      ($unsigned(wire582) ?
                          (reg588 ~^ wire569) : $unsigned(reg611)) : wire570)) : reg607[(2'h3):(2'h3)]);
              reg614 <= (~({forvar586} ?
                  ($unsigned(wire551[(3'h6):(1'h0)]) ?
                      {$unsigned(reg593),
                          wire571} : ($signed(reg612) <= (~wire549))) : reg606[(2'h3):(1'h0)]));
            end
          if (reg589)
            begin
              reg615 = (reg565 ^~ ($signed($signed(((8'hb3) ?
                      reg581 : reg604))) ?
                  (^$signed(wire547)) : ({$signed(forvar591), (~reg596)} ?
                      (~&$signed(wire568)) : $signed((8'hb7)))));
              reg616 = $signed($unsigned((~reg607[(1'h0):(1'h0)])));
              reg617 = reg589[(3'h6):(3'h4)];
              reg618 <= {reg587[(3'h6):(3'h4)], reg604[(1'h0):(1'h0)]};
            end
          else
            begin
              reg618 <= $unsigned({$signed((~^{reg595, reg565}))});
              reg619 = (&$unsigned({$unsigned((reg558 & reg615))}));
              reg620 = (forvar590[(3'h7):(3'h5)] ?
                  $signed($signed((~^(wire571 >>> (8'hb9))))) : reg606);
            end
        end
      for (forvar621 = (1'h0); (forvar621 < (2'h3)); forvar621 = (forvar621 + (1'h1)))
        begin
          for (forvar622 = (1'h0); (forvar622 < (3'h4)); forvar622 = (forvar622 + (1'h1)))
            begin
              reg623 <= ($unsigned($unsigned($unsigned(reg620[(3'h4):(2'h3)]))) * ($unsigned($unsigned(((8'hac) <<< wire569))) ?
                  (reg611[(4'ha):(1'h1)] ?
                      reg619[(3'h6):(3'h4)] : (reg562 ?
                          (~^reg593) : $unsigned(reg584))) : (wire554[(1'h0):(1'h0)] >> {(reg611 | (7'h43))})));
              reg624 = ($signed((($signed(forvar609) ?
                          (reg610 - reg606) : reg607[(3'h4):(3'h4)]) ?
                      reg587[(3'h7):(3'h6)] : forvar591[(3'h7):(2'h2)])) ?
                  reg594[(4'h8):(4'h8)] : $signed(reg605));
              reg625 <= $unsigned(((($signed(wire549) ?
                      $unsigned((8'ha6)) : (reg602 | reg565)) ?
                  $signed(((8'ha2) ?
                      reg604 : reg604)) : (~wire548[(2'h3):(1'h1)])) ^~ reg619[(5'h10):(3'h5)]));
            end
        end
    end
  assign wire626 = (-(($unsigned(reg588) ?
                       ($unsigned(reg562) == (~(8'hb7))) : (-((8'hb6) ?
                           wire548 : wire555))) ^~ $signed($unsigned(reg595[(3'h4):(2'h2)]))));
  assign wire627 = {{$signed($signed((reg598 ? wire554 : reg581))),
                           (wire626 >= {((8'hb1) ? (8'h9c) : reg580)})}};
  assign wire628 = ((+(reg604 <= $unsigned($unsigned((8'ha0))))) ?
                       ($signed(((wire547 ? reg561 : wire548) || reg581)) ?
                           (reg618[(4'hc):(1'h0)] ?
                               (|reg558) : (wire555 ?
                                   $unsigned(wire566) : $signed(wire570))) : reg588) : ({$signed((^~reg608))} & $signed(((8'hae) ?
                           wire549 : (wire548 ? wire555 : (8'ha8))))));
  assign wire629 = $signed($signed((reg594 >>> ($signed(wire571) ?
                       $unsigned(wire568) : $signed(reg601)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module463  (y, clk, wire468, wire467, wire466, wire465, wire464);
  output wire [(32'h33a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire468;
  input wire signed [(5'h10):(1'h0)] wire467;
  input wire signed [(5'h14):(1'h0)] wire466;
  input wire [(4'hf):(1'h0)] wire465;
  input wire [(4'hc):(1'h0)] wire464;
  wire [(5'h15):(1'h0)] wire542;
  wire signed [(3'h5):(1'h0)] wire541;
  wire [(4'hc):(1'h0)] wire540;
  wire signed [(2'h2):(1'h0)] wire539;
  wire signed [(5'h12):(1'h0)] wire538;
  wire signed [(4'h9):(1'h0)] wire537;
  wire signed [(4'ha):(1'h0)] wire536;
  wire signed [(3'h4):(1'h0)] wire535;
  wire [(3'h6):(1'h0)] wire534;
  wire signed [(4'he):(1'h0)] wire533;
  wire [(4'hc):(1'h0)] wire532;
  wire signed [(4'ha):(1'h0)] wire472;
  wire [(2'h2):(1'h0)] wire471;
  wire [(4'h9):(1'h0)] wire470;
  wire signed [(4'hd):(1'h0)] wire469;
  reg [(5'h11):(1'h0)] reg531 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg530 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg527 = (1'h0);
  reg [(4'hb):(1'h0)] reg524 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg522 = (1'h0);
  reg [(4'hd):(1'h0)] reg521 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg520 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg519 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg518 = (1'h0);
  reg [(4'hd):(1'h0)] reg516 = (1'h0);
  reg [(4'h9):(1'h0)] reg515 = (1'h0);
  reg [(4'hb):(1'h0)] reg511 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg509 = (1'h0);
  reg [(3'h7):(1'h0)] reg508 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg504 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg494 = (1'h0);
  reg [(4'hb):(1'h0)] reg489 = (1'h0);
  reg [(3'h4):(1'h0)] reg499 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg496 = (1'h0);
  reg [(4'hd):(1'h0)] reg495 = (1'h0);
  reg [(3'h5):(1'h0)] reg493 = (1'h0);
  reg [(4'h9):(1'h0)] reg491 = (1'h0);
  reg [(4'hf):(1'h0)] reg490 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg487 = (1'h0);
  reg [(4'hb):(1'h0)] reg483 = (1'h0);
  reg [(5'h11):(1'h0)] reg482 = (1'h0);
  reg [(4'h8):(1'h0)] reg481 = (1'h0);
  reg [(4'hb):(1'h0)] reg480 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg477 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg474 = (1'h0);
  reg [(4'he):(1'h0)] reg529 = (1'h0);
  reg [(3'h6):(1'h0)] reg528 = (1'h0);
  reg [(5'h11):(1'h0)] forvar526 = (1'h0);
  reg [(4'ha):(1'h0)] reg525 = (1'h0);
  reg [(5'h11):(1'h0)] forvar523 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar517 = (1'h0);
  reg [(4'hf):(1'h0)] reg514 = (1'h0);
  reg [(4'h8):(1'h0)] forvar513 = (1'h0);
  reg [(4'he):(1'h0)] reg512 = (1'h0);
  reg [(4'h9):(1'h0)] reg510 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar507 = (1'h0);
  reg [(5'h12):(1'h0)] reg506 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg505 = (1'h0);
  reg [(4'hd):(1'h0)] forvar503 = (1'h0);
  reg [(3'h5):(1'h0)] forvar502 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar488 = (1'h0);
  reg [(4'h8):(1'h0)] reg501 = (1'h0);
  reg [(4'ha):(1'h0)] reg500 = (1'h0);
  reg [(4'h8):(1'h0)] forvar498 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg497 = (1'h0);
  reg [(5'h15):(1'h0)] forvar494 = (1'h0);
  reg [(4'hb):(1'h0)] reg492 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar489 = (1'h0);
  reg [(5'h10):(1'h0)] reg488 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg486 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg485 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar484 = (1'h0);
  reg [(3'h7):(1'h0)] reg479 = (1'h0);
  reg signed [(4'he):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar476 = (1'h0);
  reg [(4'h8):(1'h0)] reg475 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar473 = (1'h0);
  assign y = {wire542,
                 wire541,
                 wire540,
                 wire539,
                 wire538,
                 wire537,
                 wire536,
                 wire535,
                 wire534,
                 wire533,
                 wire532,
                 wire472,
                 wire471,
                 wire470,
                 wire469,
                 reg531,
                 reg530,
                 reg527,
                 reg524,
                 reg522,
                 reg521,
                 reg520,
                 reg519,
                 reg518,
                 reg516,
                 reg515,
                 reg511,
                 reg509,
                 reg508,
                 reg504,
                 reg494,
                 reg489,
                 reg499,
                 reg496,
                 reg495,
                 reg493,
                 reg491,
                 reg490,
                 reg487,
                 reg483,
                 reg482,
                 reg481,
                 reg480,
                 reg477,
                 reg474,
                 reg529,
                 reg528,
                 forvar526,
                 reg525,
                 forvar523,
                 forvar517,
                 reg514,
                 forvar513,
                 reg512,
                 reg510,
                 forvar507,
                 reg506,
                 reg505,
                 forvar503,
                 forvar502,
                 forvar488,
                 reg501,
                 reg500,
                 forvar498,
                 reg497,
                 forvar494,
                 reg492,
                 forvar489,
                 reg488,
                 reg486,
                 reg485,
                 forvar484,
                 reg479,
                 reg478,
                 forvar476,
                 reg475,
                 forvar473,
                 (1'h0)};
  assign wire469 = ((+$unsigned(($signed(wire468) * $signed(wire464)))) ?
                       (~{(8'hb7)}) : (&$unsigned(wire468)));
  assign wire470 = {(8'ha8)};
  assign wire471 = (^~wire466);
  assign wire472 = wire464;
  always
    @(posedge clk) begin
      for (forvar473 = (1'h0); (forvar473 < (2'h3)); forvar473 = (forvar473 + (1'h1)))
        begin
          reg474 <= (~^$signed((8'hb7)));
          reg475 = $unsigned({({(|wire472)} - ({wire471, wire464} ?
                  $unsigned(wire470) : {(8'hbc)}))});
          for (forvar476 = (1'h0); (forvar476 < (2'h3)); forvar476 = (forvar476 + (1'h1)))
            begin
              reg477 <= $unsigned($signed($signed((+$signed(forvar473)))));
              reg478 = $signed($signed(({wire471} ?
                  (^(&forvar473)) : (^~((8'ha1) >>> (7'h41))))));
              reg479 = ($signed(((((8'hab) ? forvar476 : reg475) ?
                      (~wire468) : (~|wire469)) ?
                  $unsigned((~^wire472)) : (wire465 ^ reg475[(2'h2):(1'h1)]))) >>> ((~^wire465) != $unsigned((~&reg475))));
              reg480 <= wire470[(3'h5):(1'h0)];
              reg481 <= (wire472 ?
                  ((^~wire469[(3'h6):(3'h4)]) || $signed($signed($signed(reg478)))) : $unsigned((8'hb6)));
            end
          reg482 <= $signed($unsigned((~&(!(reg478 || wire471)))));
        end
      reg483 <= ({$signed(($signed(reg474) > (forvar473 <<< (8'hbd))))} <<< (($unsigned((wire467 ?
              reg477 : wire465)) * ($unsigned(wire470) ?
              forvar473[(4'ha):(1'h0)] : (reg477 ? wire471 : wire468))) ?
          (^(~^(reg482 ?
              wire465 : wire470))) : $signed(forvar473[(4'h9):(3'h7)])));
      if ($unsigned((&reg475)))
        begin
          for (forvar484 = (1'h0); (forvar484 < (2'h3)); forvar484 = (forvar484 + (1'h1)))
            begin
              reg485 = (8'hac);
              reg486 = (((reg481[(2'h2):(1'h1)] ?
                  (~&wire471[(2'h2):(1'h0)]) : $unsigned(reg485)) >> (~|$unsigned((reg478 + wire468)))) > $signed((!$unsigned(reg474))));
              reg487 <= (~reg474);
              reg488 = (^wire464[(3'h4):(3'h4)]);
            end
          for (forvar489 = (1'h0); (forvar489 < (1'h0)); forvar489 = (forvar489 + (1'h1)))
            begin
              reg490 <= ($signed($unsigned(($unsigned(forvar484) ?
                      (reg483 > wire466) : reg486[(3'h5):(2'h3)]))) ?
                  forvar484 : (&($unsigned((wire466 + reg474)) ?
                      (^(&reg481)) : ((~^reg488) ?
                          $unsigned(reg478) : (reg477 >>> reg485)))));
              reg491 <= ($unsigned((-{(reg490 ? wire470 : (8'hbc)),
                  (wire469 | wire471)})) < wire470[(2'h3):(1'h0)]);
              reg492 = reg483[(4'h9):(3'h4)];
              reg493 <= (^~$signed($signed($signed((|reg492)))));
            end
          for (forvar494 = (1'h0); (forvar494 < (1'h0)); forvar494 = (forvar494 + (1'h1)))
            begin
              reg495 <= $unsigned(((~((wire464 + forvar494) ?
                  $unsigned(reg488) : reg474[(1'h1):(1'h0)])) & (&($unsigned(wire468) != (reg487 < wire469)))));
              reg496 <= $unsigned((($unsigned(reg475) && (wire464[(4'hb):(4'h9)] ?
                  (forvar494 ?
                      (8'ha3) : reg490) : $unsigned(forvar484))) || (((wire466 ?
                      forvar484 : forvar494) ?
                  (wire470 ?
                      reg485 : reg485) : {(8'ha1)}) >> ($signed((8'ha3)) == (|(8'hac))))));
              reg497 = ((|reg490[(4'hb):(2'h2)]) ?
                  $unsigned($unsigned(wire472[(4'ha):(3'h5)])) : $unsigned($signed(forvar476[(4'h8):(3'h5)])));
            end
          for (forvar498 = (1'h0); (forvar498 < (3'h4)); forvar498 = (forvar498 + (1'h1)))
            begin
              reg499 <= (8'ha7);
              reg500 = (reg474 ?
                  (8'hbd) : $signed($signed(reg481[(2'h2):(1'h0)])));
            end
          reg501 = wire464;
        end
      else
        begin
          for (forvar484 = (1'h0); (forvar484 < (3'h4)); forvar484 = (forvar484 + (1'h1)))
            begin
              reg487 <= {$signed(({{reg482}} ?
                      $unsigned($signed(reg483)) : ((forvar473 ?
                          reg482 : reg491) | (wire464 ? reg479 : reg488)))),
                  $signed($signed({(wire466 + reg483)}))};
            end
          for (forvar488 = (1'h0); (forvar488 < (2'h2)); forvar488 = (forvar488 + (1'h1)))
            begin
              reg489 <= (+((reg475 ?
                      forvar473 : {(reg481 << (8'hab)), (-reg501)}) ?
                  {reg479} : reg481));
              reg492 = $signed((forvar489 && {($signed(forvar484) ?
                      (+(8'hab)) : (reg497 ^ forvar484))}));
              reg493 <= {$signed({((^reg497) ? $unsigned(reg492) : forvar498),
                      ($signed(forvar484) < ((7'h43) >= reg486))})};
              reg494 <= reg496[(3'h5):(2'h2)];
              reg495 <= ({$unsigned({{(8'hb5)}})} << $unsigned((~|wire467[(4'hf):(4'h8)])));
            end
        end
      for (forvar502 = (1'h0); (forvar502 < (2'h3)); forvar502 = (forvar502 + (1'h1)))
        begin
          for (forvar503 = (1'h0); (forvar503 < (2'h3)); forvar503 = (forvar503 + (1'h1)))
            begin
              reg504 <= $signed((8'ha2));
              reg505 = $signed($unsigned(reg496[(2'h2):(1'h0)]));
              reg506 = wire464;
            end
          for (forvar507 = (1'h0); (forvar507 < (2'h2)); forvar507 = (forvar507 + (1'h1)))
            begin
              reg508 <= $unsigned($signed($signed((reg493 + $signed((8'hb1))))));
              reg509 <= (8'hac);
              reg510 = {($unsigned(($unsigned(forvar476) ?
                          $signed(reg504) : (wire471 ? forvar473 : (8'hae)))) ?
                      (|reg488) : ($signed(((8'h9e) ~^ reg501)) ?
                          ($signed(forvar494) <= wire470) : $unsigned($signed(wire471))))};
              reg511 <= $unsigned($unsigned($signed($unsigned({reg505}))));
            end
          reg512 = (~$signed($unsigned((reg504 * wire468))));
          for (forvar513 = (1'h0); (forvar513 < (3'h4)); forvar513 = (forvar513 + (1'h1)))
            begin
              reg514 = {($signed(reg474) ?
                      reg485 : $signed(({reg491, wire467} && (reg474 ?
                          reg478 : reg497)))),
                  ($signed(forvar488) ?
                      $unsigned(reg497) : reg477[(1'h0):(1'h0)])};
              reg515 <= (8'ha5);
              reg516 <= $signed(({forvar507[(2'h2):(1'h1)],
                      {reg487, ((8'hac) <= wire469)}} ?
                  reg500[(3'h7):(3'h4)] : $unsigned($unsigned((reg480 ?
                      wire469 : wire467)))));
            end
          for (forvar517 = (1'h0); (forvar517 < (2'h3)); forvar517 = (forvar517 + (1'h1)))
            begin
              reg518 <= ($signed(reg508) ?
                  ((wire469 ?
                          (~&reg474[(2'h2):(2'h2)]) : reg489[(2'h2):(2'h2)]) ?
                      reg478 : ($signed((!wire465)) ~^ $unsigned(forvar494[(5'h14):(5'h10)]))) : ($unsigned(reg488) >= $unsigned((~(reg516 ~^ wire467)))));
              reg519 <= forvar513;
              reg520 <= (8'hbe);
              reg521 <= ($unsigned(($signed((~^reg518)) == $unsigned($signed(reg474)))) >= (reg520 ?
                  $unsigned(reg514[(3'h5):(2'h3)]) : {reg486,
                      $unsigned((forvar489 ~^ reg491))}));
              reg522 <= ((~|$signed(reg482[(1'h0):(1'h0)])) >= $unsigned((-reg495[(4'hc):(3'h6)])));
            end
        end
      for (forvar523 = (1'h0); (forvar523 < (1'h1)); forvar523 = (forvar523 + (1'h1)))
        begin
          if (reg501[(3'h4):(2'h3)])
            begin
              reg524 <= wire467;
            end
          else
            begin
              reg525 = (forvar523[(4'ha):(1'h1)] ?
                  $signed($signed((forvar473 ?
                      forvar494[(5'h13):(4'ha)] : reg496))) : forvar507[(3'h5):(2'h3)]);
            end
          for (forvar526 = (1'h0); (forvar526 < (2'h3)); forvar526 = (forvar526 + (1'h1)))
            begin
              reg527 <= $signed(($unsigned({$unsigned(forvar489),
                  $signed(reg500)}) > ((~forvar513) ?
                  {(forvar488 || forvar526)} : reg481[(2'h2):(2'h2)])));
              reg528 = $unsigned((~^(+$unsigned(((8'haf) ?
                  reg527 : forvar502)))));
              reg529 = ((reg485 ?
                      $signed(reg477) : (~^((reg479 ?
                          reg482 : (8'haf)) & (forvar489 & wire472)))) ?
                  (8'hb9) : ($unsigned(($signed(forvar503) & $signed(reg485))) >> (($unsigned(reg506) <= (reg475 ?
                      (8'hb9) : reg520)) >= $signed(reg516))));
              reg530 <= ((reg504 ^ $unsigned((+(-wire466)))) >= reg490[(4'hd):(2'h2)]);
              reg531 <= ($unsigned(reg495[(1'h0):(1'h0)]) * (|((reg529 < $unsigned(reg492)) << ((^~reg528) ^~ $unsigned((8'hbe))))));
            end
        end
    end
  assign wire532 = wire469[(3'h7):(3'h6)];
  assign wire533 = $signed($signed(reg482[(4'hf):(4'hd)]));
  assign wire534 = $unsigned(wire469);
  assign wire535 = {{reg524[(4'ha):(2'h3)], reg491}};
  assign wire536 = $unsigned(({$signed(reg516)} <<< $unsigned(wire465[(2'h3):(2'h2)])));
  assign wire537 = ($signed((~^$unsigned((wire532 ?
                       reg508 : wire471)))) + $signed($signed({wire472,
                       (reg480 | wire533)})));
  assign wire538 = reg494;
  assign wire539 = {{{(~^(wire536 ? (8'hb6) : wire471))},
                           ({$unsigned(reg520), wire537} << $signed({wire469,
                               (8'ha0)}))},
                       $signed($unsigned(reg477[(2'h2):(2'h2)]))};
  assign wire540 = (reg518[(3'h5):(1'h1)] ?
                       $unsigned((((wire471 > reg527) >>> $signed(reg527)) ?
                           wire468[(1'h0):(1'h0)] : ((^~wire464) != (~^reg527)))) : $unsigned({(|$unsigned((8'ha9)))}));
  assign wire541 = $unsigned($signed(($signed(reg477) ?
                       ($unsigned(wire471) ?
                           (reg494 ? wire534 : reg495) : (reg490 ?
                               wire540 : reg477)) : ($signed(wire464) + (reg494 ^~ wire540)))));
  assign wire542 = (reg482 ?
                       reg509[(4'hb):(3'h7)] : (reg522 < (~(+$unsigned((8'hbf))))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module374
#(parameter param458 = ((~{((^(8'hb9)) ? ((8'ha8) ? (8'hb8) : (8'hb6)) : ((8'hac) | (8'ha0)))}) ? ((-({(8'hb4)} ? {(8'ha8), (7'h42)} : ((8'ha1) << (8'ha0)))) << (&(7'h40))) : {(((~^(8'ha4)) | (+(8'hb1))) ^ ({(7'h43), (8'ha3)} ? {(8'ha1), (8'h9e)} : ((8'hb4) ? (7'h42) : (8'hb7)))), (&(~&((8'ha5) != (8'hb8))))}), 
parameter param459 = ((~^((^(8'ha7)) ^~ (param458 && (|param458)))) ? (({{param458}, {param458, param458}} <= param458) ? (((~&param458) ? (param458 ? param458 : param458) : {param458}) ? {param458} : (param458 ~^ param458)) : ({(~^param458), param458} ? ((7'h43) | {param458}) : {(param458 ? param458 : param458)})) : ({((param458 ? param458 : param458) > (&param458)), (-(param458 >> param458))} ^ param458)))
(y, clk, wire378, wire377, wire376, wire375);
  output wire [(32'h3a6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire378;
  input wire [(4'he):(1'h0)] wire377;
  input wire [(5'h14):(1'h0)] wire376;
  input wire signed [(2'h3):(1'h0)] wire375;
  wire signed [(4'hd):(1'h0)] wire457;
  wire [(4'h9):(1'h0)] wire456;
  wire [(5'h10):(1'h0)] wire455;
  wire [(5'h12):(1'h0)] wire435;
  wire [(3'h5):(1'h0)] wire434;
  wire [(4'hf):(1'h0)] wire433;
  wire signed [(4'he):(1'h0)] wire432;
  wire signed [(4'he):(1'h0)] wire431;
  wire signed [(4'hd):(1'h0)] wire430;
  wire [(5'h12):(1'h0)] wire382;
  wire signed [(5'h15):(1'h0)] wire381;
  wire signed [(4'hc):(1'h0)] wire380;
  wire signed [(4'h8):(1'h0)] wire379;
  reg signed [(2'h2):(1'h0)] reg453 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg451 = (1'h0);
  reg [(3'h5):(1'h0)] reg448 = (1'h0);
  reg [(2'h3):(1'h0)] reg446 = (1'h0);
  reg [(4'hf):(1'h0)] reg445 = (1'h0);
  reg [(3'h4):(1'h0)] reg443 = (1'h0);
  reg [(4'hf):(1'h0)] reg439 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg438 = (1'h0);
  reg [(4'hc):(1'h0)] reg429 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg428 = (1'h0);
  reg [(5'h14):(1'h0)] reg427 = (1'h0);
  reg [(4'hb):(1'h0)] reg426 = (1'h0);
  reg [(5'h14):(1'h0)] reg424 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg423 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg417 = (1'h0);
  reg [(5'h13):(1'h0)] reg416 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg415 = (1'h0);
  reg [(4'ha):(1'h0)] reg412 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg411 = (1'h0);
  reg [(2'h2):(1'h0)] reg410 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg408 = (1'h0);
  reg [(4'hb):(1'h0)] reg400 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg399 = (1'h0);
  reg [(4'hf):(1'h0)] reg395 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg394 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg393 = (1'h0);
  reg [(4'hd):(1'h0)] reg389 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg387 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg386 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg452 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg450 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar449 = (1'h0);
  reg [(4'hb):(1'h0)] reg447 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg444 = (1'h0);
  reg [(4'ha):(1'h0)] forvar442 = (1'h0);
  reg [(4'h8):(1'h0)] reg441 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg440 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar437 = (1'h0);
  reg [(4'hb):(1'h0)] forvar436 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar425 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg422 = (1'h0);
  reg [(5'h15):(1'h0)] forvar421 = (1'h0);
  reg [(3'h4):(1'h0)] reg420 = (1'h0);
  reg [(4'hb):(1'h0)] reg419 = (1'h0);
  reg [(5'h13):(1'h0)] reg418 = (1'h0);
  reg [(3'h4):(1'h0)] forvar414 = (1'h0);
  reg [(2'h2):(1'h0)] forvar413 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar409 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg407 = (1'h0);
  reg [(5'h10):(1'h0)] reg406 = (1'h0);
  reg [(5'h11):(1'h0)] reg405 = (1'h0);
  reg [(5'h12):(1'h0)] forvar404 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg403 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar402 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg401 = (1'h0);
  reg [(3'h5):(1'h0)] reg398 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar397 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar396 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg392 = (1'h0);
  reg [(4'he):(1'h0)] reg391 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar390 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg388 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar385 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg384 = (1'h0);
  reg [(4'he):(1'h0)] forvar383 = (1'h0);
  assign y = {wire457,
                 wire456,
                 wire455,
                 wire435,
                 wire434,
                 wire433,
                 wire432,
                 wire431,
                 wire430,
                 wire382,
                 wire381,
                 wire380,
                 wire379,
                 reg453,
                 reg451,
                 reg448,
                 reg446,
                 reg445,
                 reg443,
                 reg439,
                 reg438,
                 reg429,
                 reg428,
                 reg427,
                 reg426,
                 reg424,
                 reg423,
                 reg417,
                 reg416,
                 reg415,
                 reg412,
                 reg411,
                 reg410,
                 reg408,
                 reg400,
                 reg399,
                 reg395,
                 reg394,
                 reg393,
                 reg389,
                 reg387,
                 reg386,
                 reg454,
                 reg452,
                 reg450,
                 forvar449,
                 reg447,
                 reg444,
                 forvar442,
                 reg441,
                 reg440,
                 forvar437,
                 forvar436,
                 forvar425,
                 reg422,
                 forvar421,
                 reg420,
                 reg419,
                 reg418,
                 forvar414,
                 forvar413,
                 forvar409,
                 reg407,
                 reg406,
                 reg405,
                 forvar404,
                 reg403,
                 forvar402,
                 reg401,
                 reg398,
                 forvar397,
                 forvar396,
                 reg392,
                 reg391,
                 forvar390,
                 reg388,
                 forvar385,
                 reg384,
                 forvar383,
                 (1'h0)};
  assign wire379 = wire375[(2'h3):(1'h1)];
  assign wire380 = $unsigned((|wire377));
  assign wire381 = $unsigned((&$unsigned(($signed(wire376) ?
                       (wire378 & wire378) : $signed(wire377)))));
  assign wire382 = (~|wire379);
  always
    @(posedge clk) begin
      for (forvar383 = (1'h0); (forvar383 < (1'h0)); forvar383 = (forvar383 + (1'h1)))
        begin
          reg384 = (&$unsigned($unsigned({$unsigned(wire379), (^wire380)})));
          for (forvar385 = (1'h0); (forvar385 < (2'h2)); forvar385 = (forvar385 + (1'h1)))
            begin
              reg386 <= ((($signed($signed(wire382)) ?
                          wire377[(4'h8):(4'h8)] : $unsigned($signed(wire380))) ?
                      (wire377[(3'h4):(2'h2)] == forvar385) : wire376[(3'h5):(1'h0)]) ?
                  wire381[(3'h5):(1'h1)] : forvar383);
              reg387 <= wire381[(2'h3):(2'h2)];
              reg388 = $signed($unsigned((wire380 ?
                  (~(~|wire378)) : (wire382 ?
                      $unsigned(wire379) : (+wire380)))));
              reg389 <= {($unsigned((8'ha5)) < $signed({{wire378, forvar385},
                      (+(8'ha0))})),
                  reg388[(3'h5):(2'h3)]};
            end
          for (forvar390 = (1'h0); (forvar390 < (1'h0)); forvar390 = (forvar390 + (1'h1)))
            begin
              reg391 = $signed(({(~|forvar383[(3'h4):(3'h4)])} ?
                  reg387 : wire375[(1'h1):(1'h0)]));
              reg392 = ((^{(|wire376), wire380[(1'h1):(1'h1)]}) ?
                  (~|($signed((wire382 ?
                      wire379 : wire375)) <= $unsigned((wire375 ?
                      wire382 : (8'h9c))))) : {(wire381 + $signed((wire382 >> wire375)))});
              reg393 <= forvar385[(5'h11):(4'hd)];
              reg394 <= $signed((wire378[(3'h7):(3'h5)] ?
                  (({reg388} ? reg391 : ((8'hbf) >= wire377)) ^~ ((wire381 ?
                      reg387 : reg393) >>> $unsigned(wire375))) : $signed((7'h43))));
              reg395 <= $unsigned({wire381[(3'h6):(1'h1)],
                  ($unsigned($signed(reg394)) ?
                      {forvar383} : (^~(reg386 ? reg389 : reg384)))});
            end
        end
      for (forvar396 = (1'h0); (forvar396 < (1'h0)); forvar396 = (forvar396 + (1'h1)))
        begin
          for (forvar397 = (1'h0); (forvar397 < (2'h2)); forvar397 = (forvar397 + (1'h1)))
            begin
              reg398 = $unsigned((wire375 ?
                  wire375[(1'h1):(1'h0)] : reg395[(2'h2):(1'h0)]));
              reg399 <= $unsigned((~&($unsigned(wire378[(4'h9):(1'h0)]) ?
                  reg388[(3'h5):(1'h1)] : (^~(reg391 < reg393)))));
              reg400 <= ((~$signed($unsigned((forvar397 - forvar390)))) ?
                  (|{(&reg384),
                      ((8'hbb) ?
                          $unsigned(reg398) : $signed(reg388))}) : reg394[(3'h7):(1'h1)]);
              reg401 = wire380;
            end
          for (forvar402 = (1'h0); (forvar402 < (2'h3)); forvar402 = (forvar402 + (1'h1)))
            begin
              reg403 = (!{$unsigned(wire381)});
            end
          for (forvar404 = (1'h0); (forvar404 < (2'h2)); forvar404 = (forvar404 + (1'h1)))
            begin
              reg405 = {(($signed($signed(wire378)) ?
                          $signed((~^wire380)) : $signed($signed(wire380))) ?
                      $signed(wire379[(3'h5):(2'h3)]) : ($signed(wire378[(2'h3):(2'h2)]) ?
                          {(!reg394)} : forvar390[(2'h2):(1'h1)])),
                  $unsigned($signed((~reg389[(3'h6):(3'h4)])))};
              reg406 = (($signed(((forvar383 <<< reg395) ?
                      $signed(forvar383) : (~&wire376))) ?
                  (8'had) : $signed(reg391[(4'he):(4'hd)])) ~^ $unsigned((({wire375,
                          wire377} ?
                      forvar396[(2'h2):(1'h0)] : ((8'hbb) ?
                          reg405 : forvar397)) ?
                  (forvar404[(1'h1):(1'h0)] > reg392) : $signed($unsigned(reg391)))));
              reg407 = wire376[(4'hb):(1'h0)];
              reg408 <= $unsigned((reg394[(1'h1):(1'h1)] ?
                  $unsigned($signed((reg388 ?
                      forvar390 : reg391))) : forvar396[(4'h9):(4'h9)]));
            end
          for (forvar409 = (1'h0); (forvar409 < (3'h4)); forvar409 = (forvar409 + (1'h1)))
            begin
              reg410 <= (reg408[(2'h2):(1'h1)] ?
                  ($unsigned(((reg407 || wire380) ?
                      (^forvar390) : $unsigned(wire376))) >>> reg386) : ($signed($unsigned((^wire379))) >= $unsigned((^~(wire382 ?
                      (8'hb9) : forvar402)))));
            end
        end
      reg411 <= ((-{reg394[(3'h7):(1'h0)], forvar402[(2'h2):(2'h2)]}) ?
          {$unsigned($signed((~|reg388)))} : (~^$unsigned((reg399 && (&reg386)))));
      reg412 <= (~^(!$signed(($signed((7'h42)) ?
          (forvar396 || reg403) : reg393))));
      for (forvar413 = (1'h0); (forvar413 < (1'h0)); forvar413 = (forvar413 + (1'h1)))
        begin
          for (forvar414 = (1'h0); (forvar414 < (1'h1)); forvar414 = (forvar414 + (1'h1)))
            begin
              reg415 <= (reg399 + ((+reg406) * (($signed(wire379) >= $signed(reg395)) ^ ((~^forvar409) & reg403))));
              reg416 <= $signed($unsigned((reg415 ?
                  ((wire379 ?
                      wire381 : wire376) < $signed(reg387)) : ((+reg386) || $signed(reg412)))));
              reg417 <= $signed((^~$unsigned(($unsigned(reg395) ?
                  $unsigned(reg401) : forvar385[(4'he):(4'h9)]))));
              reg418 = ($signed({{$unsigned(wire377)}}) + (8'ha5));
              reg419 = (~|$unsigned(reg398[(3'h5):(2'h3)]));
            end
          reg420 = (~&reg410);
          for (forvar421 = (1'h0); (forvar421 < (1'h0)); forvar421 = (forvar421 + (1'h1)))
            begin
              reg422 = (&reg419[(3'h5):(3'h4)]);
              reg423 <= reg399[(4'hb):(3'h7)];
              reg424 <= reg410[(2'h2):(2'h2)];
            end
          for (forvar425 = (1'h0); (forvar425 < (2'h3)); forvar425 = (forvar425 + (1'h1)))
            begin
              reg426 <= ($unsigned((~|(~forvar409))) << {reg419[(2'h3):(2'h2)]});
              reg427 <= forvar383;
              reg428 <= $unsigned($unsigned(((&(^reg423)) + {$unsigned(forvar425)})));
            end
          reg429 <= (($unsigned((reg386 | $signed((8'ha1)))) ?
                  (8'hb7) : wire378) ?
              $signed((($signed((8'hb6)) ?
                      $unsigned(forvar396) : $signed(reg418)) ?
                  (-reg420[(3'h4):(1'h1)]) : reg416[(4'he):(4'ha)])) : reg419[(4'h8):(1'h0)]);
        end
    end
  assign wire430 = $unsigned({$unsigned((reg429[(4'h8):(3'h6)] ?
                           (8'h9f) : reg393[(5'h10):(3'h6)])),
                       (-($unsigned(wire378) ?
                           (wire379 ~^ wire380) : (-reg417)))});
  assign wire431 = reg394[(2'h2):(1'h0)];
  assign wire432 = wire380[(1'h1):(1'h0)];
  assign wire433 = (8'h9f);
  assign wire434 = $unsigned($signed({wire377}));
  assign wire435 = $signed($signed($signed({reg429[(1'h0):(1'h0)],
                       (reg394 && reg394)})));
  always
    @(posedge clk) begin
      for (forvar436 = (1'h0); (forvar436 < (2'h2)); forvar436 = (forvar436 + (1'h1)))
        begin
          for (forvar437 = (1'h0); (forvar437 < (1'h0)); forvar437 = (forvar437 + (1'h1)))
            begin
              reg438 <= reg412[(3'h6):(3'h6)];
              reg439 <= (-$unsigned(wire430));
              reg440 = reg389;
            end
          reg441 = (!reg394);
          for (forvar442 = (1'h0); (forvar442 < (2'h3)); forvar442 = (forvar442 + (1'h1)))
            begin
              reg443 <= reg387;
              reg444 = (reg394[(3'h7):(1'h1)] ?
                  ((forvar436 ?
                          ((-reg441) >>> (reg415 * (8'hbf))) : ((reg394 ?
                                  wire435 : reg441) ?
                              (~^wire379) : $unsigned(reg415))) ?
                      wire376[(2'h2):(1'h1)] : (7'h43)) : reg416);
              reg445 <= (((-reg444) >>> reg423) ?
                  (((reg410 ? (reg438 ? (8'hbe) : reg410) : $unsigned(reg412)) ?
                          (-(-reg410)) : (^~reg408)) ?
                      ((~|(~wire377)) ?
                          ((wire430 >= wire430) <<< wire435) : {$unsigned(reg410)}) : (+$signed($signed(reg387)))) : (reg439[(4'h9):(4'h9)] ~^ ((^$unsigned(reg428)) ?
                      $signed($unsigned((8'ha9))) : ((+reg440) < (wire432 && (8'hb0))))));
              reg446 <= $unsigned((~^reg412));
              reg447 = ((-reg441[(3'h6):(2'h3)]) << $signed(reg416[(2'h3):(1'h0)]));
            end
          reg448 <= $signed($unsigned(((wire378[(2'h3):(2'h3)] <<< forvar442) ?
              forvar436 : (-wire377[(2'h2):(1'h1)]))));
          for (forvar449 = (1'h0); (forvar449 < (3'h4)); forvar449 = (forvar449 + (1'h1)))
            begin
              reg450 = $unsigned({$unsigned($signed($signed(reg393)))});
              reg451 <= wire430[(4'hc):(2'h2)];
              reg452 = $unsigned(forvar442);
              reg453 <= {{(+wire380[(3'h7):(2'h2)])}};
            end
        end
      reg454 = ((wire381[(4'h8):(3'h6)] ?
              $signed($signed(reg393[(4'hf):(4'h9)])) : reg452) ?
          reg441 : $unsigned($unsigned((reg452[(1'h0):(1'h0)] + {(8'hbf)}))));
    end
  assign wire455 = reg438;
  assign wire456 = reg427[(4'hb):(4'h8)];
  assign wire457 = ($signed(reg439[(3'h4):(2'h3)]) != (({(-(8'haf)),
                               {(7'h42)}} ?
                           wire430 : (wire377[(4'h9):(4'h9)] ?
                               (+wire433) : (+(7'h44)))) ?
                       $signed($unsigned($signed((8'hab)))) : $signed($signed(((8'ha2) <= reg424)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module292
#(parameter param370 = (~((8'ha1) - ((((7'h42) ? (8'ha0) : (8'hb4)) ? ((8'h9e) ? (8'ha8) : (7'h42)) : (~&(8'hb3))) * (((8'ha8) ? (8'ha2) : (8'h9c)) ? (8'ha5) : ((8'haa) ? (8'hb0) : (8'ha8)))))), 
parameter param371 = (8'hb2))
(y, clk, wire296, wire295, wire294, wire293);
  output wire [(32'h372):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire296;
  input wire signed [(3'h6):(1'h0)] wire295;
  input wire signed [(5'h14):(1'h0)] wire294;
  input wire [(5'h15):(1'h0)] wire293;
  wire signed [(4'hb):(1'h0)] wire369;
  wire signed [(4'hf):(1'h0)] wire368;
  wire signed [(4'hd):(1'h0)] wire367;
  wire [(5'h10):(1'h0)] wire366;
  wire signed [(5'h13):(1'h0)] wire365;
  wire [(5'h12):(1'h0)] wire364;
  wire signed [(3'h5):(1'h0)] wire363;
  wire signed [(5'h11):(1'h0)] wire362;
  wire [(4'hb):(1'h0)] wire361;
  wire [(4'ha):(1'h0)] wire360;
  wire signed [(2'h2):(1'h0)] wire359;
  wire signed [(4'hb):(1'h0)] wire358;
  wire signed [(5'h15):(1'h0)] wire357;
  wire signed [(4'h8):(1'h0)] wire356;
  wire [(5'h10):(1'h0)] wire355;
  wire [(4'he):(1'h0)] wire354;
  wire signed [(5'h15):(1'h0)] wire353;
  wire [(5'h10):(1'h0)] wire352;
  wire [(4'hd):(1'h0)] wire351;
  wire signed [(4'hf):(1'h0)] wire350;
  wire [(3'h6):(1'h0)] wire297;
  reg signed [(4'ha):(1'h0)] reg347 = (1'h0);
  reg [(4'hd):(1'h0)] reg345 = (1'h0);
  reg [(4'hb):(1'h0)] reg344 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg341 = (1'h0);
  reg [(5'h13):(1'h0)] reg338 = (1'h0);
  reg [(4'h8):(1'h0)] reg337 = (1'h0);
  reg [(4'hb):(1'h0)] reg332 = (1'h0);
  reg [(5'h10):(1'h0)] reg331 = (1'h0);
  reg [(5'h14):(1'h0)] reg327 = (1'h0);
  reg [(4'hf):(1'h0)] reg324 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg322 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg321 = (1'h0);
  reg [(3'h4):(1'h0)] reg319 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg318 = (1'h0);
  reg [(5'h11):(1'h0)] reg317 = (1'h0);
  reg signed [(4'he):(1'h0)] reg316 = (1'h0);
  reg signed [(4'he):(1'h0)] reg314 = (1'h0);
  reg [(4'hd):(1'h0)] reg311 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg310 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg309 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg307 = (1'h0);
  reg [(5'h11):(1'h0)] reg306 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg303 = (1'h0);
  reg [(5'h14):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg300 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg349 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg348 = (1'h0);
  reg [(3'h4):(1'h0)] reg346 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar343 = (1'h0);
  reg [(5'h13):(1'h0)] reg342 = (1'h0);
  reg [(4'he):(1'h0)] forvar340 = (1'h0);
  reg [(4'hb):(1'h0)] forvar339 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar336 = (1'h0);
  reg [(4'hd):(1'h0)] reg335 = (1'h0);
  reg [(4'he):(1'h0)] reg334 = (1'h0);
  reg [(3'h7):(1'h0)] forvar333 = (1'h0);
  reg [(5'h13):(1'h0)] reg330 = (1'h0);
  reg [(4'h9):(1'h0)] forvar329 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg328 = (1'h0);
  reg [(2'h3):(1'h0)] forvar326 = (1'h0);
  reg [(4'hc):(1'h0)] forvar325 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg323 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar320 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar315 = (1'h0);
  reg [(4'h8):(1'h0)] forvar313 = (1'h0);
  reg [(2'h3):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar308 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar305 = (1'h0);
  reg [(3'h5):(1'h0)] forvar304 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg301 = (1'h0);
  reg [(5'h15):(1'h0)] forvar299 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar298 = (1'h0);
  assign y = {wire369,
                 wire368,
                 wire367,
                 wire366,
                 wire365,
                 wire364,
                 wire363,
                 wire362,
                 wire361,
                 wire360,
                 wire359,
                 wire358,
                 wire357,
                 wire356,
                 wire355,
                 wire354,
                 wire353,
                 wire352,
                 wire351,
                 wire350,
                 wire297,
                 reg347,
                 reg345,
                 reg344,
                 reg341,
                 reg338,
                 reg337,
                 reg332,
                 reg331,
                 reg327,
                 reg324,
                 reg322,
                 reg321,
                 reg319,
                 reg318,
                 reg317,
                 reg316,
                 reg314,
                 reg311,
                 reg310,
                 reg309,
                 reg307,
                 reg306,
                 reg303,
                 reg302,
                 reg300,
                 reg349,
                 reg348,
                 reg346,
                 forvar343,
                 reg342,
                 forvar340,
                 forvar339,
                 forvar336,
                 reg335,
                 reg334,
                 forvar333,
                 reg330,
                 forvar329,
                 reg328,
                 forvar326,
                 forvar325,
                 reg323,
                 forvar320,
                 forvar315,
                 forvar313,
                 reg312,
                 forvar308,
                 forvar305,
                 forvar304,
                 reg301,
                 forvar299,
                 forvar298,
                 (1'h0)};
  assign wire297 = (!(wire294[(4'hc):(2'h3)] ?
                       ($signed((wire296 + (8'hbf))) > wire295) : (($unsigned(wire294) ?
                           (wire295 ?
                               wire295 : wire296) : $signed(wire293)) != wire294)));
  always
    @(posedge clk) begin
      for (forvar298 = (1'h0); (forvar298 < (3'h4)); forvar298 = (forvar298 + (1'h1)))
        begin
          for (forvar299 = (1'h0); (forvar299 < (2'h2)); forvar299 = (forvar299 + (1'h1)))
            begin
              reg300 <= wire296;
              reg301 = $signed((($signed((~wire293)) && $signed($unsigned((8'hb0)))) ?
                  (((forvar298 ?
                      wire297 : forvar299) != (-wire294)) != $unsigned($signed(wire294))) : (forvar299 - (8'hb8))));
              reg302 <= $unsigned(forvar298);
              reg303 <= {reg302, (wire293 << ($signed(wire293) | reg300))};
            end
        end
      for (forvar304 = (1'h0); (forvar304 < (1'h0)); forvar304 = (forvar304 + (1'h1)))
        begin
          for (forvar305 = (1'h0); (forvar305 < (1'h1)); forvar305 = (forvar305 + (1'h1)))
            begin
              reg306 <= $unsigned(wire297[(3'h6):(2'h2)]);
              reg307 <= reg301;
            end
          for (forvar308 = (1'h0); (forvar308 < (1'h0)); forvar308 = (forvar308 + (1'h1)))
            begin
              reg309 <= $unsigned(reg301);
              reg310 <= $unsigned(wire296);
              reg311 <= $signed($signed($signed((|(wire296 ?
                  wire296 : wire295)))));
              reg312 = $unsigned(((($unsigned(reg300) ?
                  (forvar304 ?
                      (8'hb2) : forvar308) : reg302) || forvar308) | $signed(($unsigned(wire294) ?
                  forvar298 : (~|(8'ha2))))));
            end
          for (forvar313 = (1'h0); (forvar313 < (1'h1)); forvar313 = (forvar313 + (1'h1)))
            begin
              reg314 <= reg309;
            end
          for (forvar315 = (1'h0); (forvar315 < (1'h0)); forvar315 = (forvar315 + (1'h1)))
            begin
              reg316 <= ((~|$unsigned($unsigned($unsigned(reg306)))) ~^ $signed(($unsigned($unsigned((7'h41))) ?
                  ((wire293 ?
                      (8'ha2) : (8'ha7)) <<< reg312[(2'h2):(2'h2)]) : reg307[(2'h3):(1'h0)])));
              reg317 <= $signed((((!$signed((8'ha0))) ?
                      forvar308 : ((~^forvar298) ? $signed(wire296) : reg310)) ?
                  reg316[(2'h3):(1'h1)] : ((((7'h43) != forvar313) || (reg310 ?
                      forvar298 : forvar298)) * $unsigned((^~reg303)))));
              reg318 <= $unsigned(forvar305[(1'h0):(1'h0)]);
              reg319 <= reg302;
            end
          for (forvar320 = (1'h0); (forvar320 < (2'h2)); forvar320 = (forvar320 + (1'h1)))
            begin
              reg321 <= (^{$signed($signed((^forvar305))),
                  ({(7'h42),
                      $signed(reg318)} << $unsigned(reg309[(1'h0):(1'h0)]))});
              reg322 <= {$unsigned((~^wire297[(2'h2):(1'h1)])),
                  forvar315[(4'hd):(3'h7)]};
              reg323 = reg319;
              reg324 <= (($unsigned((~|(forvar298 ? reg323 : reg307))) ?
                      $signed((reg318 ^~ forvar305)) : (forvar320[(1'h0):(1'h0)] >>> ($unsigned(reg321) ^~ reg310[(1'h1):(1'h0)]))) ?
                  $signed($unsigned(reg309[(4'hd):(4'h8)])) : reg322[(3'h5):(2'h3)]);
            end
        end
      for (forvar325 = (1'h0); (forvar325 < (1'h1)); forvar325 = (forvar325 + (1'h1)))
        begin
          for (forvar326 = (1'h0); (forvar326 < (3'h4)); forvar326 = (forvar326 + (1'h1)))
            begin
              reg327 <= (reg300[(4'hd):(2'h2)] >> (-forvar305));
              reg328 = (+(~&(&{(reg314 ? reg302 : forvar304), reg327})));
            end
          for (forvar329 = (1'h0); (forvar329 < (1'h0)); forvar329 = (forvar329 + (1'h1)))
            begin
              reg330 = $signed($unsigned(($signed(wire293) ?
                  (^$signed(reg309)) : (wire295 ?
                      (forvar329 ? (8'hb9) : reg301) : (reg306 ?
                          reg314 : forvar329)))));
              reg331 <= (((forvar329 ?
                      (reg328[(2'h3):(2'h3)] ?
                          (~forvar320) : $unsigned(forvar298)) : ($unsigned(reg321) ?
                          (forvar326 ? reg309 : reg324) : $unsigned((7'h40)))) ?
                  $unsigned(reg309[(3'h6):(2'h3)]) : (|(^~$unsigned(wire293)))) ~^ {$unsigned((forvar315[(4'hf):(4'h9)] | forvar320[(2'h2):(1'h0)])),
                  reg310[(3'h6):(1'h1)]});
              reg332 <= wire297[(3'h4):(3'h4)];
            end
          for (forvar333 = (1'h0); (forvar333 < (1'h1)); forvar333 = (forvar333 + (1'h1)))
            begin
              reg334 = reg307;
              reg335 = (~|reg301);
            end
          for (forvar336 = (1'h0); (forvar336 < (3'h4)); forvar336 = (forvar336 + (1'h1)))
            begin
              reg337 <= (-wire293[(4'hb):(4'h9)]);
              reg338 <= reg309[(4'hc):(2'h3)];
            end
        end
      for (forvar339 = (1'h0); (forvar339 < (1'h1)); forvar339 = (forvar339 + (1'h1)))
        begin
          for (forvar340 = (1'h0); (forvar340 < (2'h2)); forvar340 = (forvar340 + (1'h1)))
            begin
              reg341 <= (8'hb0);
            end
          reg342 = forvar304[(2'h2):(2'h2)];
          for (forvar343 = (1'h0); (forvar343 < (2'h3)); forvar343 = (forvar343 + (1'h1)))
            begin
              reg344 <= forvar339;
            end
          if (($signed($signed($unsigned((reg306 ? forvar305 : forvar308)))) ?
              $unsigned((((forvar299 ? reg310 : reg307) ?
                      forvar299[(5'h11):(4'hf)] : $signed(reg317)) ?
                  forvar340 : ($signed(wire296) ^ reg301[(2'h2):(1'h1)]))) : forvar340))
            begin
              reg345 <= ((-reg317[(3'h4):(1'h0)]) ?
                  reg317[(4'hc):(3'h7)] : reg334);
              reg346 = (($signed($unsigned((reg310 ^ reg317))) ^~ reg330[(3'h5):(2'h2)]) ?
                  $unsigned(((forvar333 ?
                      $signed(forvar298) : (!forvar333)) << forvar298)) : (^$unsigned(reg318[(2'h3):(1'h0)])));
              reg347 <= $signed(((^((forvar313 - (8'ha1)) ?
                      $signed((7'h42)) : $unsigned((8'hba)))) ?
                  {((reg307 ?
                          (8'h9f) : (8'hb0)) ~^ (+(8'ha8)))} : {$unsigned($unsigned(reg300))}));
            end
          else
            begin
              reg346 = (($unsigned(reg342[(1'h1):(1'h0)]) ?
                      reg317[(1'h1):(1'h0)] : $signed((wire294[(4'ha):(2'h3)] ?
                          $signed(reg316) : {reg332}))) ?
                  (reg334[(1'h0):(1'h0)] | {reg303[(3'h4):(3'h4)],
                      forvar339}) : $unsigned(forvar298));
              reg347 <= reg322[(2'h2):(1'h1)];
              reg348 = (~&(({wire297,
                  $unsigned(forvar304)} << (forvar343 | (wire297 == reg323))) ~^ $unsigned(forvar305)));
            end
        end
      reg349 = (^((^~$unsigned($unsigned((8'h9e)))) + ($unsigned(forvar315) ?
          (((8'hbc) < reg335) == (forvar304 == (7'h43))) : reg323[(2'h2):(2'h2)])));
    end
  assign wire350 = (8'ha8);
  assign wire351 = (~^reg310);
  assign wire352 = ((~|wire294[(5'h14):(2'h2)]) | reg309);
  assign wire353 = reg309[(4'h9):(1'h0)];
  assign wire354 = ({(~(~^(reg319 ?
                           reg318 : reg331)))} & reg317[(4'he):(4'he)]);
  assign wire355 = reg310[(1'h1):(1'h0)];
  assign wire356 = (8'hb1);
  assign wire357 = (8'hbd);
  assign wire358 = ($signed({(reg314 >= (reg306 ? reg322 : reg302)),
                           $unsigned((reg319 && reg331))}) ?
                       $signed($unsigned((wire293[(2'h2):(1'h0)] & (reg306 ?
                           reg341 : reg314)))) : wire354);
  assign wire359 = wire355;
  assign wire360 = reg302;
  assign wire361 = $unsigned(((7'h43) ~^ (!$unsigned({reg300}))));
  assign wire362 = $unsigned($unsigned(wire359));
  assign wire363 = ($signed(reg302[(5'h11):(4'hb)]) > (&$signed((-(~|reg322)))));
  assign wire364 = reg344[(4'ha):(3'h4)];
  assign wire365 = $unsigned((((&$unsigned(reg347)) ?
                       $unsigned($signed(reg331)) : $unsigned($unsigned(reg306))) >= ($signed((^~reg345)) ?
                       wire353 : $unsigned((reg311 ? wire353 : reg318)))));
  assign wire366 = $unsigned($signed(reg331));
  assign wire367 = (({($signed((8'h9c)) <<< $unsigned(reg306)),
                           (wire365[(5'h10):(2'h2)] << (wire293 ^ wire294))} ^~ ($unsigned((reg311 ?
                               wire353 : wire355)) ?
                           ((reg337 < (8'ha1)) - wire360[(1'h0):(1'h0)]) : $unsigned($unsigned(wire358)))) ?
                       $unsigned(($unsigned((!wire356)) >> (|$signed((8'had))))) : (^$unsigned(((wire294 <<< wire361) ?
                           wire365 : (~wire353)))));
  assign wire368 = $unsigned($signed(((((8'ha4) == (8'hac)) ?
                           (reg309 < reg300) : (8'hba)) ?
                       $unsigned({wire356}) : ((+reg302) ~^ {wire294}))));
  assign wire369 = (~|$unsigned($unsigned(reg327)));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module167  (y, clk, wire171, wire170, wire169, wire168);
  output wire [(32'h4de):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire171;
  input wire [(3'h4):(1'h0)] wire170;
  input wire signed [(4'ha):(1'h0)] wire169;
  input wire [(4'he):(1'h0)] wire168;
  wire [(5'h10):(1'h0)] wire289;
  wire [(4'hd):(1'h0)] wire288;
  wire signed [(3'h7):(1'h0)] wire287;
  wire [(4'he):(1'h0)] wire244;
  wire signed [(4'ha):(1'h0)] wire243;
  wire [(2'h2):(1'h0)] wire242;
  wire [(4'hb):(1'h0)] wire204;
  wire signed [(5'h12):(1'h0)] wire172;
  reg signed [(3'h7):(1'h0)] reg286 = (1'h0);
  reg [(4'hc):(1'h0)] reg284 = (1'h0);
  reg [(4'hd):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg278 = (1'h0);
  reg [(5'h13):(1'h0)] reg274 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg273 = (1'h0);
  reg signed [(4'he):(1'h0)] reg272 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg271 = (1'h0);
  reg [(3'h7):(1'h0)] reg268 = (1'h0);
  reg [(4'hd):(1'h0)] reg267 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg266 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg265 = (1'h0);
  reg [(2'h2):(1'h0)] reg262 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg261 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg260 = (1'h0);
  reg [(4'he):(1'h0)] reg257 = (1'h0);
  reg [(4'ha):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg255 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg254 = (1'h0);
  reg [(4'h8):(1'h0)] reg253 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg250 = (1'h0);
  reg [(4'hf):(1'h0)] reg248 = (1'h0);
  reg [(4'h9):(1'h0)] reg247 = (1'h0);
  reg [(4'hb):(1'h0)] reg238 = (1'h0);
  reg [(2'h2):(1'h0)] reg237 = (1'h0);
  reg [(4'hf):(1'h0)] reg235 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg228 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg225 = (1'h0);
  reg [(4'he):(1'h0)] reg221 = (1'h0);
  reg [(3'h5):(1'h0)] reg220 = (1'h0);
  reg [(5'h10):(1'h0)] reg219 = (1'h0);
  reg [(4'hf):(1'h0)] reg216 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg215 = (1'h0);
  reg [(3'h5):(1'h0)] reg212 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg210 = (1'h0);
  reg [(2'h3):(1'h0)] reg209 = (1'h0);
  reg [(3'h4):(1'h0)] reg203 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg202 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg201 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg200 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg198 = (1'h0);
  reg [(4'hd):(1'h0)] reg196 = (1'h0);
  reg [(4'hc):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg189 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg188 = (1'h0);
  reg [(4'hf):(1'h0)] reg186 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg184 = (1'h0);
  reg [(4'h9):(1'h0)] reg183 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg181 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg180 = (1'h0);
  reg [(4'hb):(1'h0)] reg178 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg177 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg176 = (1'h0);
  reg [(4'hf):(1'h0)] reg285 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar283 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar282 = (1'h0);
  reg [(5'h12):(1'h0)] reg281 = (1'h0);
  reg [(3'h6):(1'h0)] reg280 = (1'h0);
  reg [(2'h2):(1'h0)] reg277 = (1'h0);
  reg [(4'hb):(1'h0)] forvar276 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg275 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar270 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar269 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar264 = (1'h0);
  reg [(4'hd):(1'h0)] reg263 = (1'h0);
  reg [(4'he):(1'h0)] forvar259 = (1'h0);
  reg [(2'h2):(1'h0)] forvar258 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg252 = (1'h0);
  reg [(4'ha):(1'h0)] forvar251 = (1'h0);
  reg [(3'h4):(1'h0)] reg249 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar246 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar245 = (1'h0);
  reg [(3'h6):(1'h0)] reg241 = (1'h0);
  reg [(5'h11):(1'h0)] reg240 = (1'h0);
  reg [(4'he):(1'h0)] reg239 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar236 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar234 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar233 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg231 = (1'h0);
  reg [(4'h8):(1'h0)] forvar230 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar227 = (1'h0);
  reg [(3'h4):(1'h0)] forvar226 = (1'h0);
  reg [(4'hc):(1'h0)] forvar224 = (1'h0);
  reg [(5'h14):(1'h0)] reg223 = (1'h0);
  reg [(4'hd):(1'h0)] forvar222 = (1'h0);
  reg [(2'h2):(1'h0)] forvar218 = (1'h0);
  reg [(2'h3):(1'h0)] forvar217 = (1'h0);
  reg [(5'h12):(1'h0)] forvar214 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg213 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg211 = (1'h0);
  reg [(5'h10):(1'h0)] reg208 = (1'h0);
  reg [(2'h2):(1'h0)] forvar207 = (1'h0);
  reg [(4'he):(1'h0)] reg206 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar205 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg199 = (1'h0);
  reg [(2'h2):(1'h0)] forvar197 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg195 = (1'h0);
  reg [(4'h8):(1'h0)] forvar194 = (1'h0);
  reg [(5'h13):(1'h0)] forvar193 = (1'h0);
  reg [(5'h14):(1'h0)] reg192 = (1'h0);
  reg [(5'h12):(1'h0)] reg190 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar187 = (1'h0);
  reg [(4'he):(1'h0)] forvar185 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg182 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar175 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg174 = (1'h0);
  reg [(4'he):(1'h0)] forvar173 = (1'h0);
  assign y = {wire289,
                 wire288,
                 wire287,
                 wire244,
                 wire243,
                 wire242,
                 wire204,
                 wire172,
                 reg286,
                 reg284,
                 reg279,
                 reg278,
                 reg274,
                 reg273,
                 reg272,
                 reg271,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg262,
                 reg261,
                 reg260,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg253,
                 reg250,
                 reg248,
                 reg247,
                 reg238,
                 reg237,
                 reg235,
                 reg232,
                 reg228,
                 reg225,
                 reg221,
                 reg220,
                 reg219,
                 reg216,
                 reg215,
                 reg212,
                 reg210,
                 reg209,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg198,
                 reg196,
                 reg191,
                 reg189,
                 reg188,
                 reg186,
                 reg184,
                 reg183,
                 reg181,
                 reg180,
                 reg178,
                 reg177,
                 reg176,
                 reg285,
                 forvar283,
                 forvar282,
                 reg281,
                 reg280,
                 reg277,
                 forvar276,
                 reg275,
                 forvar270,
                 forvar269,
                 forvar264,
                 reg263,
                 forvar259,
                 forvar258,
                 reg252,
                 forvar251,
                 reg249,
                 forvar246,
                 forvar245,
                 reg241,
                 reg240,
                 reg239,
                 forvar236,
                 forvar234,
                 forvar233,
                 reg231,
                 forvar230,
                 reg229,
                 forvar227,
                 forvar226,
                 forvar224,
                 reg223,
                 forvar222,
                 forvar218,
                 forvar217,
                 forvar214,
                 reg213,
                 reg211,
                 reg208,
                 forvar207,
                 reg206,
                 forvar205,
                 reg199,
                 forvar197,
                 reg195,
                 forvar194,
                 forvar193,
                 reg192,
                 reg190,
                 forvar187,
                 forvar185,
                 reg182,
                 reg179,
                 forvar175,
                 reg174,
                 forvar173,
                 (1'h0)};
  assign wire172 = ($signed(($signed($signed((8'h9d))) ?
                       ($signed(wire168) < (wire171 ?
                           wire171 : wire169)) : $unsigned(wire170[(2'h3):(1'h0)]))) - $signed((wire170[(1'h1):(1'h1)] ?
                       wire170 : (wire170 >> (8'had)))));
  always
    @(posedge clk) begin
      for (forvar173 = (1'h0); (forvar173 < (3'h4)); forvar173 = (forvar173 + (1'h1)))
        begin
          reg174 = (~^((^~(wire171[(3'h4):(1'h1)] ?
                  ((8'hb2) ? wire170 : wire172) : (wire172 ?
                      wire168 : wire172))) ?
              wire170 : $signed((~(wire172 ? wire172 : (8'haf))))));
          for (forvar175 = (1'h0); (forvar175 < (2'h3)); forvar175 = (forvar175 + (1'h1)))
            begin
              reg176 <= (({(wire168[(4'ha):(2'h3)] ?
                              $unsigned(forvar173) : (forvar175 ?
                                  forvar173 : (7'h40)))} ?
                      (^~((forvar173 ?
                          wire171 : forvar173) == $unsigned(wire172))) : wire171[(4'hd):(4'hc)]) ?
                  (+(wire169 & $signed($unsigned(wire168)))) : forvar175[(4'hf):(3'h5)]);
              reg177 <= $signed((((^wire171) ?
                      $unsigned((!forvar173)) : reg174[(4'h9):(3'h6)]) ?
                  $unsigned(forvar173) : wire170[(2'h2):(1'h0)]));
              reg178 <= $signed(((!$unsigned((!wire168))) << wire172[(4'hd):(2'h3)]));
              reg179 = ((^~$signed(forvar175)) ?
                  $signed($unsigned({$signed(reg178)})) : $unsigned($signed((forvar175[(1'h1):(1'h1)] << (wire171 ?
                      (7'h42) : forvar173)))));
              reg180 <= $unsigned($signed($unsigned($unsigned((8'h9c)))));
            end
          if ((&$unsigned((reg178[(4'h9):(4'h9)] ?
              $signed((wire171 ? wire171 : wire168)) : reg179))))
            begin
              reg181 <= ((~$signed({reg180, (8'h9e)})) ?
                  (-reg174[(4'ha):(3'h7)]) : $signed($unsigned($unsigned({wire168}))));
              reg182 = $unsigned(wire171);
            end
          else
            begin
              reg181 <= (!(reg178[(3'h6):(3'h5)] ^ (~&$unsigned($unsigned(wire170)))));
              reg183 <= ({(~&(reg178[(2'h3):(1'h1)] - reg176)),
                  reg181} < (((~((8'ha9) ? forvar175 : reg174)) & {(~wire170),
                      (~^(8'h9f))}) ?
                  reg180 : (~wire168)));
              reg184 <= $signed($unsigned(reg179));
            end
          for (forvar185 = (1'h0); (forvar185 < (1'h0)); forvar185 = (forvar185 + (1'h1)))
            begin
              reg186 <= ((~^(~&$signed(reg182))) ?
                  ({(+$unsigned(reg182))} ^ reg180[(2'h3):(1'h1)]) : forvar185);
            end
          for (forvar187 = (1'h0); (forvar187 < (3'h4)); forvar187 = (forvar187 + (1'h1)))
            begin
              reg188 <= reg176[(3'h6):(2'h3)];
              reg189 <= reg181;
              reg190 = (((reg176 && $unsigned($signed(forvar185))) ^~ $signed(((^~wire172) ?
                      $signed(forvar185) : {(8'hb8), forvar187}))) ?
                  (wire169 && $unsigned(({reg186} ?
                      $unsigned(reg179) : $unsigned((7'h43))))) : $signed(reg179));
              reg191 <= (~(forvar187[(3'h7):(3'h7)] ?
                  (^~((~&reg180) ?
                      wire168[(3'h5):(1'h1)] : (forvar187 ?
                          reg174 : reg188))) : $signed(wire171[(4'he):(4'hb)])));
            end
        end
      reg192 = (($unsigned(((8'hb5) ?
              (~|reg176) : (reg180 < (8'hbe)))) >> forvar175[(4'hd):(1'h0)]) ?
          reg174[(3'h6):(3'h4)] : {$unsigned({(reg184 ? forvar175 : forvar173),
                  $signed((8'hb4))}),
              (reg182[(1'h1):(1'h1)] ?
                  (forvar185[(1'h1):(1'h1)] ?
                      {reg178} : (reg182 == reg183)) : $signed({reg190,
                      reg177}))});
      for (forvar193 = (1'h0); (forvar193 < (1'h0)); forvar193 = (forvar193 + (1'h1)))
        begin
          for (forvar194 = (1'h0); (forvar194 < (3'h4)); forvar194 = (forvar194 + (1'h1)))
            begin
              reg195 = reg181[(4'h9):(2'h3)];
              reg196 <= ($signed(reg183) <= (~(&reg190)));
            end
          for (forvar197 = (1'h0); (forvar197 < (1'h0)); forvar197 = (forvar197 + (1'h1)))
            begin
              reg198 <= ($signed(((~((8'hb1) ? reg192 : reg182)) ?
                      {$unsigned((8'ha5)), (reg181 > reg174)} : {(reg176 ?
                              (8'hb7) : forvar197),
                          {reg182, forvar193}})) ?
                  (^reg188[(1'h1):(1'h0)]) : (forvar185[(2'h2):(1'h0)] ?
                      reg190[(4'hc):(4'ha)] : wire170));
              reg199 = wire171;
              reg200 <= {(~|{((forvar194 ?
                          reg189 : wire170) < $signed(reg177))}),
                  forvar197};
            end
          reg201 <= ((~|$signed(((&forvar175) > forvar187))) < ((^~(+(reg182 ?
                  forvar197 : reg190))) ?
              ((~^$unsigned(reg180)) ?
                  reg199[(4'hb):(4'ha)] : (~&(reg190 ?
                      reg191 : forvar185))) : {(!reg184[(3'h5):(1'h1)])}));
          reg202 <= reg199[(4'h9):(1'h0)];
          reg203 <= $signed(((!((8'hb7) ? reg186 : (&reg178))) ?
              $signed($unsigned((~^forvar173))) : reg184[(4'ha):(1'h1)]));
        end
    end
  assign wire204 = (|reg198);
  always
    @(posedge clk) begin
      for (forvar205 = (1'h0); (forvar205 < (1'h1)); forvar205 = (forvar205 + (1'h1)))
        begin
          reg206 = wire170;
          for (forvar207 = (1'h0); (forvar207 < (1'h1)); forvar207 = (forvar207 + (1'h1)))
            begin
              reg208 = ({$signed((reg201 ~^ $unsigned(reg203))),
                      (!((reg181 ? wire169 : wire169) >>> $signed(reg198)))} ?
                  wire170 : reg191);
              reg209 <= {$unsigned(({(reg183 & reg201), wire171} ?
                      reg176 : $unsigned(reg181))),
                  (reg206 - $signed((^reg203)))};
              reg210 <= ((&$signed(reg177)) ?
                  $signed((~$unsigned(reg178))) : $signed(($signed((reg191 & (8'ha9))) ?
                      (^(reg181 > reg177)) : $signed(reg181))));
              reg211 = $signed($unsigned(wire172[(5'h12):(4'h8)]));
              reg212 <= $signed(wire168[(1'h0):(1'h0)]);
            end
          reg213 = $signed(reg183[(3'h4):(1'h0)]);
          for (forvar214 = (1'h0); (forvar214 < (2'h2)); forvar214 = (forvar214 + (1'h1)))
            begin
              reg215 <= reg203;
              reg216 <= (-{$signed($signed($unsigned(reg212)))});
            end
        end
      for (forvar217 = (1'h0); (forvar217 < (2'h2)); forvar217 = (forvar217 + (1'h1)))
        begin
          for (forvar218 = (1'h0); (forvar218 < (1'h0)); forvar218 = (forvar218 + (1'h1)))
            begin
              reg219 <= (~^$unsigned((-$signed((reg198 * (8'haf))))));
              reg220 <= reg184[(1'h1):(1'h0)];
            end
          reg221 <= (!$signed(($unsigned(((7'h40) & reg220)) ?
              $unsigned(reg200) : ((reg183 == forvar205) ?
                  (!(8'hae)) : $signed(reg213)))));
          for (forvar222 = (1'h0); (forvar222 < (1'h0)); forvar222 = (forvar222 + (1'h1)))
            begin
              reg223 = (^~($unsigned($signed(reg186)) != $signed((&reg196))));
            end
          for (forvar224 = (1'h0); (forvar224 < (2'h2)); forvar224 = (forvar224 + (1'h1)))
            begin
              reg225 <= ({$signed((8'had))} <= (^~$unsigned(({reg188} ~^ $signed(reg203)))));
            end
        end
      for (forvar226 = (1'h0); (forvar226 < (3'h4)); forvar226 = (forvar226 + (1'h1)))
        begin
          for (forvar227 = (1'h0); (forvar227 < (1'h0)); forvar227 = (forvar227 + (1'h1)))
            begin
              reg228 <= (-{(-((8'hb2) ? forvar224 : $signed(reg176))),
                  reg188[(1'h1):(1'h0)]});
              reg229 = $unsigned(forvar217);
            end
          for (forvar230 = (1'h0); (forvar230 < (1'h0)); forvar230 = (forvar230 + (1'h1)))
            begin
              reg231 = $unsigned($signed($unsigned(((forvar226 ?
                  (8'hbd) : forvar217) || (~|forvar230)))));
            end
          reg232 <= ((~reg177) || $signed(((reg213 ?
                  $unsigned(forvar207) : (forvar218 ? reg228 : forvar224)) ?
              reg189 : ((reg208 << reg213) ? {reg184} : (wire171 >> reg216)))));
        end
      for (forvar233 = (1'h0); (forvar233 < (2'h3)); forvar233 = (forvar233 + (1'h1)))
        begin
          for (forvar234 = (1'h0); (forvar234 < (1'h1)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 <= (|{$signed((&reg181[(3'h4):(2'h2)]))});
            end
          for (forvar236 = (1'h0); (forvar236 < (3'h4)); forvar236 = (forvar236 + (1'h1)))
            begin
              reg237 <= ((reg201 >= ({$signed(reg200),
                  forvar236} + $signed($unsigned(forvar214)))) ^~ (wire170 <= ((-(~|reg201)) && reg180)));
              reg238 <= ($unsigned($signed(forvar234)) >> reg178);
              reg239 = wire172[(3'h4):(2'h2)];
              reg240 = (~^((~|$signed((reg186 - reg238))) | $unsigned($unsigned(forvar230))));
              reg241 = (wire204[(2'h3):(2'h2)] >> $unsigned($unsigned(($signed((8'hb5)) == (8'ha6)))));
            end
        end
    end
  assign wire242 = (^(~({reg203[(2'h3):(1'h0)], {reg183, reg209}} && reg200)));
  assign wire243 = (reg209[(1'h1):(1'h1)] ?
                       $signed(reg176[(2'h2):(1'h1)]) : (^~wire242[(1'h0):(1'h0)]));
  assign wire244 = $signed((~wire243[(4'ha):(3'h5)]));
  always
    @(posedge clk) begin
      for (forvar245 = (1'h0); (forvar245 < (2'h2)); forvar245 = (forvar245 + (1'h1)))
        begin
          for (forvar246 = (1'h0); (forvar246 < (2'h3)); forvar246 = (forvar246 + (1'h1)))
            begin
              reg247 <= reg235[(2'h2):(2'h2)];
              reg248 <= reg232;
              reg249 = {wire243[(3'h5):(2'h3)], wire172[(4'h8):(4'h8)]};
              reg250 <= $unsigned(reg180);
            end
          for (forvar251 = (1'h0); (forvar251 < (3'h4)); forvar251 = (forvar251 + (1'h1)))
            begin
              reg252 = reg200;
              reg253 <= ((reg203 > forvar251[(4'ha):(3'h7)]) ~^ reg200[(4'h8):(3'h6)]);
              reg254 <= (reg247[(3'h6):(1'h1)] | $signed(reg198));
            end
          reg255 <= ((~&((reg198[(4'h9):(3'h5)] ?
                  reg247[(3'h7):(3'h6)] : (^~reg249)) ?
              $signed($unsigned(reg184)) : (reg216 ?
                  reg235[(2'h2):(1'h1)] : (reg176 ?
                      reg184 : (8'ha8))))) ^~ (($unsigned($unsigned(reg235)) >>> reg216) - {reg219[(1'h1):(1'h1)]}));
          reg256 <= {(($unsigned($unsigned(wire168)) <= ($unsigned(reg184) <<< (8'hb0))) ?
                  $unsigned((~|reg249)) : reg235[(4'hf):(3'h6)]),
              reg220[(1'h1):(1'h0)]};
          reg257 <= (~|{reg176});
        end
      for (forvar258 = (1'h0); (forvar258 < (1'h0)); forvar258 = (forvar258 + (1'h1)))
        begin
          for (forvar259 = (1'h0); (forvar259 < (2'h2)); forvar259 = (forvar259 + (1'h1)))
            begin
              reg260 <= (!(-reg201[(2'h2):(1'h1)]));
              reg261 <= reg180;
              reg262 <= wire171;
              reg263 = (^(~^(reg247 ?
                  reg178 : $unsigned(wire168[(4'hd):(2'h3)]))));
            end
          for (forvar264 = (1'h0); (forvar264 < (1'h0)); forvar264 = (forvar264 + (1'h1)))
            begin
              reg265 <= reg262[(2'h2):(2'h2)];
              reg266 <= ((^reg181[(4'h9):(3'h6)]) * (|reg203));
              reg267 <= reg181[(3'h4):(2'h3)];
              reg268 <= $signed(($unsigned(reg212[(1'h0):(1'h0)]) ?
                  $signed(reg188) : ((+reg221) & forvar245)));
            end
        end
      for (forvar269 = (1'h0); (forvar269 < (2'h3)); forvar269 = (forvar269 + (1'h1)))
        begin
          for (forvar270 = (1'h0); (forvar270 < (1'h1)); forvar270 = (forvar270 + (1'h1)))
            begin
              reg271 <= (reg221 >> wire243[(3'h4):(2'h2)]);
            end
          reg272 <= reg178[(3'h5):(1'h0)];
          reg273 <= {($signed(reg200) ?
                  {(+$signed((8'hab)))} : ($signed(reg228[(3'h7):(1'h1)]) ?
                      {(reg215 <<< (8'hbe))} : ((reg249 < reg272) ?
                          (reg232 >= wire244) : $signed(wire171)))),
              reg178};
          reg274 <= $signed((^reg237[(1'h1):(1'h1)]));
          reg275 = {($unsigned(reg184) ?
                  $signed((8'ha7)) : ($signed((reg180 ? (8'hb8) : wire171)) ?
                      $signed(reg250) : forvar246)),
              forvar245[(3'h4):(2'h2)]};
        end
      for (forvar276 = (1'h0); (forvar276 < (2'h3)); forvar276 = (forvar276 + (1'h1)))
        begin
          if ((((8'hb6) >>> (reg203 * $signed((reg201 > reg228)))) ?
              $unsigned($unsigned(wire170)) : (((reg273[(3'h4):(3'h4)] ?
                      (reg250 ? reg252 : (8'ha9)) : (wire204 ?
                          reg176 : reg274)) ?
                  ((8'hb6) < (forvar276 ?
                      (8'ha3) : wire244)) : ((wire168 < reg272) ?
                      reg201[(1'h1):(1'h0)] : (reg228 ?
                          wire172 : forvar251))) != $unsigned((reg180 ?
                  $signed((8'ha0)) : (^~reg198))))))
            begin
              reg277 = (+$signed((^~(~(8'hbe)))));
            end
          else
            begin
              reg278 <= $unsigned((8'ha7));
              reg279 <= $unsigned(($signed(wire170[(2'h2):(1'h1)]) || (-reg176[(1'h0):(1'h0)])));
              reg280 = reg235[(3'h4):(1'h1)];
              reg281 = ((({(forvar270 ? wire172 : (8'ha6))} ?
                      (~(^~reg176)) : $signed((|(8'hae)))) >> reg274[(3'h4):(1'h1)]) ?
                  ((^~$signed($unsigned(reg220))) ?
                      $signed($signed($unsigned(reg216))) : $unsigned(reg272[(4'h8):(1'h0)])) : reg272[(4'hd):(4'h8)]);
            end
        end
      for (forvar282 = (1'h0); (forvar282 < (1'h1)); forvar282 = (forvar282 + (1'h1)))
        begin
          for (forvar283 = (1'h0); (forvar283 < (2'h3)); forvar283 = (forvar283 + (1'h1)))
            begin
              reg284 <= reg216;
              reg285 = reg202[(3'h4):(3'h4)];
            end
          reg286 <= (~^(forvar245 << reg202[(4'h8):(3'h4)]));
        end
    end
  assign wire287 = ($signed((8'hbf)) >= reg267);
  assign wire288 = {{reg250}};
  assign wire289 = (|(|{wire171[(4'he):(4'hd)], wire242[(2'h2):(1'h1)]}));
endmodule