(* use_dsp48="no" *) (* use_dsp="no" *) module top
#( parameter param695 = {{(8'ha9), (~&(+((7'h44) && (8'ha7))))}, (-(-(~&((8'hac) ? (7'h48) : (8'ha4)))))} )
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h295):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire0;
  input wire signed [(2'h3):(1'h0)] wire1;
  input wire [(4'hf):(1'h0)] wire2;
  input wire signed [(5'h14):(1'h0)] wire3;
  input wire signed [(4'hf):(1'h0)] wire4;
  wire [(4'hc):(1'h0)] wire694;
  wire [(5'h12):(1'h0)] wire693;
  wire [(4'h9):(1'h0)] wire692;
  wire signed [(5'h17):(1'h0)] wire691;
  wire signed [(5'h11):(1'h0)] wire690;
  reg [(3'h6):(1'h0)] forvar5 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar6 = (1'h0);
  reg [(5'h16):(1'h0)] reg7 = (1'h0);
  reg signed [(4'he):(1'h0)] reg8 = (1'h0);
  reg [(4'h8):(1'h0)] reg9 = (1'h0);
  reg [(5'h13):(1'h0)] forvar10 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg12 = (1'h0);
  reg [(3'h7):(1'h0)] reg13 = (1'h0);
  reg [(4'hb):(1'h0)] forvar14 = (1'h0);
  reg [(5'h11):(1'h0)] reg15 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg17 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg18 = (1'h0);
  reg [(5'h16):(1'h0)] reg19 = (1'h0);
  reg [(3'h7):(1'h0)] reg20 = (1'h0);
  reg [(5'h14):(1'h0)] reg21 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg22 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg23 = (1'h0);
  reg [(5'h15):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg25 = (1'h0);
  reg [(3'h6):(1'h0)] reg26 = (1'h0);
  reg [(4'hc):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg28 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg29 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg30 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg31 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg32 = (1'h0);
  reg [(5'h14):(1'h0)] reg33 = (1'h0);
  wire [(3'h4):(1'h0)] wire34;
  wire signed [(5'h15):(1'h0)] wire677;
  wire signed [(4'he):(1'h0)] wire679;
  wire [(5'h13):(1'h0)] wire680;
  wire [(4'hb):(1'h0)] wire681;
  wire signed [(5'h16):(1'h0)] wire682;
  wire [(5'h10):(1'h0)] wire683;
  wire [(5'h14):(1'h0)] wire684;
  wire signed [(4'hb):(1'h0)] wire685;
  wire [(3'h7):(1'h0)] wire686;
  wire signed [(5'h11):(1'h0)] wire687;
  wire signed [(4'hc):(1'h0)] wire688;
  assign y = {wire694,
                 wire693,
                 wire692,
                 wire691,
                 wire690,
                 forvar5,
                 forvar6,
                 reg7,
                 reg8,
                 reg9,
                 forvar10,
                 reg11,
                 reg12,
                 reg13,
                 forvar14,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg20,
                 reg21,
                 reg22,
                 reg23,
                 reg24,
                 reg25,
                 reg26,
                 reg27,
                 reg28,
                 reg29,
                 reg30,
                 reg31,
                 reg32,
                 reg33,
                 wire34,
                 wire677,
                 wire679,
                 wire680,
                 wire681,
                 wire682,
                 wire683,
                 wire684,
                 wire685,
                 wire686,
                 wire687,
                 wire688,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar5 = (1'h0); (forvar5 < (1'h1)); forvar5 = (forvar5 + (1'h1)))
        begin
          for (forvar6 = (1'h0); (forvar6 < (1'h0)); forvar6 = (forvar6 + (1'h1)))
            begin
              reg7 <= wire1;
              reg8 <= forvar6[(4'ha):(4'ha)];
              reg9 <= (8'hb6);
            end
          for (forvar10 = (1'h0); (forvar10 < (1'h1)); forvar10 = (forvar10 + (1'h1)))
            begin
              reg11 <= $signed(forvar5);
            end
        end
      reg12 <= reg7;
      reg13 <= "TTgvoZmed9nJ9CS";
      for (forvar14 = (1'h0); (forvar14 < (3'h4)); forvar14 = (forvar14 + (1'h1)))
        begin
          reg15 <= (~|(reg8[(1'h0):(1'h0)] ^~ ((^(forvar14 ?
              forvar5 : (8'ha2))) + (reg11 ? (-forvar6) : (&(8'hbe))))));
          if ((wire4 ^~ ($unsigned((^(forvar6 ?
              wire2 : (7'h40)))) ~^ wire3[(3'h5):(1'h0)])))
            begin
              reg16 <= wire0;
              reg17 <= forvar14[(2'h3):(1'h1)];
              reg18 <= (reg13[(3'h6):(2'h2)] << forvar5);
              reg19 <= ((8'ha0) || (~|wire4));
              reg20 <= ($signed(reg16) < "oCEYI");
            end
          else
            begin
              reg16 = reg16[(3'h5):(3'h5)];
            end
          if (reg11[(4'h9):(3'h5)])
            begin
              reg21 <= (forvar6 && "KtqRlGMauiP");
            end
          else
            begin
              reg21 <= (~$signed(($unsigned((-reg18)) ?
                  ((+reg18) >> (reg17 != reg19)) : $signed(wire3[(2'h2):(1'h0)]))));
              reg22 <= (&reg11);
            end
          if (reg9[(1'h0):(1'h0)])
            begin
              reg23 <= reg15;
            end
          else
            begin
              reg23 <= ((($unsigned(reg9) ~^ wire2[(3'h7):(3'h6)]) ?
                      $signed("kdyq4KCfNu0tuWBByC") : (8'h9f)) ?
                  (~|$signed($unsigned(reg19[(5'h13):(3'h4)]))) : ((8'hb0) ?
                      reg19[(4'he):(3'h4)] : ((!wire4) == $signed($signed(wire1)))));
              reg24 <= (wire1 ~^ ($signed(("DB8PWCxisCy3cJTDwP0V" ?
                  "pHS71yYLArmBt" : $unsigned(reg19))) >= $signed(((reg17 ?
                  forvar5 : (7'h48)) || "aNoOEl4OP2I"))));
              reg25 <= {(($unsigned((+wire2)) ?
                          "rYad" : $unsigned(reg15[(4'hc):(4'h8)])) ?
                      reg15[(3'h6):(3'h5)] : wire1)};
              reg26 <= "WBQTk";
              reg27 <= (forvar5[(1'h0):(1'h0)] << (8'ha1));
            end
          if ((&{(!$signed($unsigned(reg19)))}))
            begin
              reg28 <= reg18[(1'h0):(1'h0)];
              reg29 <= {(8'ha7), reg26[(2'h3):(2'h3)]};
              reg30 = reg23;
              reg31 <= $signed($signed((~$unsigned($signed(wire0)))));
            end
          else
            begin
              reg28 <= $signed((^~$unsigned(($unsigned(reg8) ?
                  wire3[(4'hf):(3'h6)] : (reg15 || forvar6)))));
              reg29 <= $unsigned($signed(""));
              reg30 <= (!"06LnF7Pym6i1o98Wss5CQ");
              reg31 <= reg23;
              reg32 <= $unsigned(reg15[(1'h0):(1'h0)]);
            end
        end
      reg33 <= "TibAIc8ZcKox";
    end
  assign wire34 = (($unsigned($unsigned((-reg16))) <<< "FpK9xAv") ?
                      reg31 : ($unsigned("ddW87cM3MY") >= (reg31 ?
                          (^reg20) : ((reg25 ~^ reg21) ^~ "wqBDku3Ml"))));
  module35 modinst678 (.wire38(reg17), .y(wire677), .wire39(reg22), .clk(clk), .wire37(reg19), .wire36(reg29));
  assign wire679 = $unsigned(((~"vq4ieJU8uzUFv0Ka") ?
                       reg16[(1'h1):(1'h1)] : $signed(wire1[(1'h1):(1'h1)])));
  assign wire680 = "Rf";
  assign wire681 = $unsigned(forvar10[(5'h13):(4'h8)]);
  assign wire682 = wire0[(3'h4):(3'h4)];
  assign wire683 = "q1vfigtdsSl82GG";
  assign wire684 = (!{wire680,
                       $unsigned(((wire2 ? (8'hbe) : wire3) ?
                           $unsigned(wire679) : reg29[(4'ha):(2'h2)]))});
  assign wire685 = (~|reg32[(1'h1):(1'h1)]);
  assign wire686 = $signed(((!reg33) ? reg27 : {reg22, "UVIwRMznPJK4fuoORF"}));
  assign wire687 = ($signed(forvar14) ~^ (~&reg33[(1'h0):(1'h0)]));
  module200 modinst689 (.clk(clk), .y(wire688), .wire205(reg7), .wire204(wire687), .wire202(reg33), .wire201(wire4), .wire203(forvar14));
  assign wire690 = ($signed("IeB") ?
                       (forvar10 ?
                           "JRTh55KL33di643Y" : "mD9sOQqsNXoWgGSRbm86Y") : (~wire680[(5'h10):(4'h9)]));
  assign wire691 = "";
  assign wire692 = ($unsigned("ss7ibaSVwHvPCQi2qUBE") + $signed($signed($signed((wire685 >= wire683)))));
  assign wire693 = $unsigned((((wire685[(3'h7):(3'h5)] ?
                       wire685 : reg18[(2'h3):(1'h1)]) - (|"4SSmPOREQJIl")) ^~ "AoUFZwgpuit4NFbme"));
  assign wire694 = (8'ha6);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module35
#( parameter param676 = ((((~&((8'ha1) ? (8'hb1) : (8'hb5))) ? (((7'h48) ? (7'h41) : (8'ha2)) ? ((7'h47) | (7'h47)) : {(8'hb9)}) : {(+(8'ha7))}) + (((^~(8'ha2)) ? (^(8'hb2)) : ((8'ha7) ? (8'haa) : (7'h42))) ? {((7'h47) || (8'h9e))} : (((7'h42) ? (8'hbc) : (8'hb8)) ? (^~(8'ha1)) : ((7'h43) ? (8'hbf) : (8'haa))))) ? (({{(8'haa)}} ? (((7'h45) + (8'ha8)) ? ((8'hb7) <= (8'ha1)) : ((8'hbc) & (7'h42))) : ((&(8'hac)) << (&(7'h47)))) ? ((&(~|(7'h44))) - (((8'hbc) ? (7'h48) : (8'ha3)) == ((8'hb9) < (7'h42)))) : (&(!((8'hb4) == (7'h45))))) : {((|((8'ha6) != (8'haa))) > (&((8'hb6) << (8'hbe))))}) )
(y, clk, wire36, wire37, wire38, wire39);
  output wire [(32'hd6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h17):(1'h0)] wire36;
  input wire signed [(5'h14):(1'h0)] wire37;
  input wire [(4'hf):(1'h0)] wire38;
  input wire signed [(5'h16):(1'h0)] wire39;
  wire [(4'he):(1'h0)] wire675;
  wire signed [(5'h14):(1'h0)] wire674;
  wire [(4'h8):(1'h0)] wire673;
  wire [(3'h6):(1'h0)] wire672;
  wire [(5'h14):(1'h0)] wire671;
  wire [(4'hb):(1'h0)] wire670;
  wire signed [(5'h14):(1'h0)] wire669;
  wire [(2'h3):(1'h0)] wire668;
  wire [(4'he):(1'h0)] wire667;
  wire signed [(3'h7):(1'h0)] wire665;
  wire [(4'he):(1'h0)] wire664;
  wire signed [(4'h8):(1'h0)] wire663;
  wire [(5'h13):(1'h0)] wire662;
  wire [(4'hb):(1'h0)] wire660;
  wire signed [(5'h12):(1'h0)] wire40;
  wire signed [(5'h14):(1'h0)] wire658;
  assign y = {wire675,
                 wire674,
                 wire673,
                 wire672,
                 wire671,
                 wire670,
                 wire669,
                 wire668,
                 wire667,
                 wire665,
                 wire664,
                 wire663,
                 wire662,
                 wire660,
                 wire40,
                 wire658,
                 (1'h0)};
  assign wire40 = (wire38 != wire38);
  module41 modinst659 (.wire43(wire40), .wire44(wire36), .wire45(wire39), .wire46(wire38), .y(wire658), .wire42(wire37), .clk(clk));
  module313 modinst661 (wire660, clk, wire40, wire39, wire658, wire38);
  assign wire662 = ((wire658 != $signed($signed((wire658 == wire38)))) & (~^wire36));
  assign wire663 = ({wire40[(3'h5):(2'h2)],
                       {((wire39 ? wire658 : wire37) ? {wire38} : "Y"),
                           "lyU8K2zA1L"}} <= (!($signed($unsigned((8'haa))) > wire662[(4'h9):(3'h7)])));
  assign wire664 = $signed((wire40[(3'h5):(2'h2)] > $unsigned(({wire660} >> $signed(wire40)))));
  module193 modinst666 (.wire197(wire658), .wire195(wire660), .wire194(wire37), .wire196(wire39), .y(wire665), .clk(clk));
  assign wire667 = wire663[(3'h5):(3'h5)];
  assign wire668 = (~|wire38);
  assign wire669 = {wire665, $unsigned($signed({wire37}))};
  assign wire670 = "lQEkT6N93O8lmuVn";
  assign wire671 = $unsigned($unsigned($signed(wire663[(1'h1):(1'h0)])));
  assign wire672 = $signed(wire663);
  assign wire673 = wire665;
  assign wire674 = $unsigned(wire662[(5'h12):(1'h1)]);
  assign wire675 = $signed("YlSoPU5uLBrV");
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module41  (y, clk, wire46, wire45, wire44, wire43, wire42);
  output wire [(32'h929):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire46;
  input wire signed [(5'h16):(1'h0)] wire45;
  input wire signed [(5'h17):(1'h0)] wire44;
  input wire [(5'h12):(1'h0)] wire43;
  input wire signed [(5'h12):(1'h0)] wire42;
  reg signed [(5'h11):(1'h0)] reg652 = (1'h0);
  reg [(4'he):(1'h0)] forvar651 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg650 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar646 = (1'h0);
  reg [(4'h9):(1'h0)] reg657 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg656 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg655 = (1'h0);
  reg [(4'hc):(1'h0)] reg654 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg653 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar652 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg651 = (1'h0);
  reg [(5'h15):(1'h0)] forvar650 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg649 = (1'h0);
  reg [(4'hf):(1'h0)] reg648 = (1'h0);
  reg [(3'h4):(1'h0)] reg647 = (1'h0);
  reg [(5'h17):(1'h0)] reg646 = (1'h0);
  reg [(4'ha):(1'h0)] reg645 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg644 = (1'h0);
  reg [(4'hc):(1'h0)] reg643 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg642 = (1'h0);
  reg [(5'h10):(1'h0)] forvar641 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg640 = (1'h0);
  reg [(5'h12):(1'h0)] reg639 = (1'h0);
  reg [(2'h2):(1'h0)] reg638 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg637 = (1'h0);
  reg [(4'hb):(1'h0)] reg636 = (1'h0);
  reg [(5'h13):(1'h0)] reg635 = (1'h0);
  reg [(5'h15):(1'h0)] forvar634 = (1'h0);
  reg [(5'h13):(1'h0)] reg633 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar625 = (1'h0);
  reg [(4'h8):(1'h0)] reg632 = (1'h0);
  reg [(2'h2):(1'h0)] reg631 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg630 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg629 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg628 = (1'h0);
  reg [(2'h2):(1'h0)] reg627 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg626 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg623 = (1'h0);
  reg [(5'h16):(1'h0)] reg622 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg621 = (1'h0);
  reg [(5'h13):(1'h0)] forvar620 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg619 = (1'h0);
  wire [(3'h6):(1'h0)] wire618;
  reg [(5'h14):(1'h0)] reg617 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg616 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar615 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg614 = (1'h0);
  reg [(5'h11):(1'h0)] reg613 = (1'h0);
  reg [(3'h7):(1'h0)] reg612 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg611 = (1'h0);
  reg [(2'h3):(1'h0)] reg610 = (1'h0);
  reg [(4'he):(1'h0)] reg609 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg608 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg607 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar606 = (1'h0);
  reg [(5'h13):(1'h0)] reg605 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg604 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar603 = (1'h0);
  reg [(5'h15):(1'h0)] reg602 = (1'h0);
  reg [(3'h5):(1'h0)] forvar601 = (1'h0);
  reg [(4'h9):(1'h0)] reg600 = (1'h0);
  reg [(5'h14):(1'h0)] reg599 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg598 = (1'h0);
  reg [(5'h13):(1'h0)] forvar597 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar596 = (1'h0);
  reg [(5'h17):(1'h0)] reg595 = (1'h0);
  reg [(5'h12):(1'h0)] reg594 = (1'h0);
  reg [(4'ha):(1'h0)] reg593 = (1'h0);
  reg [(4'ha):(1'h0)] reg592 = (1'h0);
  reg [(3'h7):(1'h0)] reg591 = (1'h0);
  reg [(5'h10):(1'h0)] reg590 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg589 = (1'h0);
  reg [(5'h15):(1'h0)] forvar588 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg587 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg586 = (1'h0);
  reg [(4'hf):(1'h0)] reg585 = (1'h0);
  reg [(3'h5):(1'h0)] reg584 = (1'h0);
  reg [(4'he):(1'h0)] reg583 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg582 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg581 = (1'h0);
  reg [(5'h16):(1'h0)] forvar580 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg579 = (1'h0);
  reg [(2'h3):(1'h0)] reg578 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar577 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg576 = (1'h0);
  reg [(4'h8):(1'h0)] reg575 = (1'h0);
  reg [(4'h9):(1'h0)] reg574 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar573 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar572 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg571 = (1'h0);
  wire signed [(5'h12):(1'h0)] wire154;
  wire [(4'h8):(1'h0)] wire156;
  wire signed [(5'h17):(1'h0)] wire157;
  wire signed [(4'hb):(1'h0)] wire158;
  reg [(5'h17):(1'h0)] forvar159 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg160 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg161 = (1'h0);
  reg [(3'h4):(1'h0)] reg162 = (1'h0);
  reg [(5'h15):(1'h0)] reg163 = (1'h0);
  reg [(2'h2):(1'h0)] forvar164 = (1'h0);
  reg [(5'h14):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg166 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg167 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg168 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg169 = (1'h0);
  reg [(4'hd):(1'h0)] forvar170 = (1'h0);
  reg [(5'h15):(1'h0)] reg171 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg172 = (1'h0);
  reg [(4'hc):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar174 = (1'h0);
  reg [(5'h15):(1'h0)] reg175 = (1'h0);
  reg signed [(4'he):(1'h0)] reg176 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar177 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg178 = (1'h0);
  reg [(3'h4):(1'h0)] reg179 = (1'h0);
  reg [(5'h10):(1'h0)] reg180 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg181 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg182 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg183 = (1'h0);
  reg [(5'h14):(1'h0)] reg184 = (1'h0);
  reg [(4'h8):(1'h0)] reg185 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar186 = (1'h0);
  reg [(5'h17):(1'h0)] reg187 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg188 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg189 = (1'h0);
  reg [(4'ha):(1'h0)] forvar190 = (1'h0);
  reg [(4'h8):(1'h0)] reg191 = (1'h0);
  wire signed [(2'h3):(1'h0)] wire192;
  wire signed [(5'h16):(1'h0)] wire525;
  wire [(4'hd):(1'h0)] wire527;
  wire [(2'h2):(1'h0)] wire528;
  wire signed [(3'h4):(1'h0)] wire529;
  wire signed [(5'h11):(1'h0)] wire530;
  reg [(4'ha):(1'h0)] forvar531 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg532 = (1'h0);
  reg [(5'h15):(1'h0)] reg533 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg534 = (1'h0);
  reg [(5'h14):(1'h0)] reg535 = (1'h0);
  reg [(4'h9):(1'h0)] reg536 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg537 = (1'h0);
  reg [(5'h10):(1'h0)] reg538 = (1'h0);
  reg [(5'h17):(1'h0)] reg539 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg540 = (1'h0);
  reg [(5'h14):(1'h0)] reg541 = (1'h0);
  reg [(3'h4):(1'h0)] reg542 = (1'h0);
  reg [(2'h2):(1'h0)] reg543 = (1'h0);
  reg [(5'h15):(1'h0)] reg544 = (1'h0);
  reg [(4'hc):(1'h0)] reg545 = (1'h0);
  reg [(5'h11):(1'h0)] reg531 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg546 = (1'h0);
  reg [(4'h9):(1'h0)] reg547 = (1'h0);
  reg [(4'hc):(1'h0)] reg548 = (1'h0);
  reg [(5'h17):(1'h0)] reg549 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg550 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg551 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg552 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg553 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg554 = (1'h0);
  reg [(3'h7):(1'h0)] reg555 = (1'h0);
  reg [(4'hc):(1'h0)] reg556 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg557 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar548 = (1'h0);
  reg [(4'hc):(1'h0)] reg558 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar559 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg560 = (1'h0);
  reg [(5'h14):(1'h0)] reg561 = (1'h0);
  reg [(3'h4):(1'h0)] reg562 = (1'h0);
  reg [(5'h13):(1'h0)] reg563 = (1'h0);
  wire [(5'h15):(1'h0)] wire564;
  wire signed [(5'h14):(1'h0)] wire565;
  wire [(4'hc):(1'h0)] wire566;
  wire signed [(5'h17):(1'h0)] wire567;
  wire [(5'h15):(1'h0)] wire568;
  wire signed [(4'h8):(1'h0)] wire569;
  assign y = {reg652,
                 forvar651,
                 reg650,
                 forvar646,
                 reg657,
                 reg656,
                 reg655,
                 reg654,
                 reg653,
                 forvar652,
                 reg651,
                 forvar650,
                 reg649,
                 reg648,
                 reg647,
                 reg646,
                 reg645,
                 reg644,
                 reg643,
                 reg642,
                 forvar641,
                 reg640,
                 reg639,
                 reg638,
                 reg637,
                 reg636,
                 reg635,
                 forvar634,
                 reg633,
                 forvar625,
                 reg632,
                 reg631,
                 reg630,
                 reg629,
                 reg628,
                 reg627,
                 reg626,
                 reg625,
                 reg624,
                 reg623,
                 reg622,
                 reg621,
                 forvar620,
                 reg619,
                 wire618,
                 reg617,
                 reg616,
                 forvar615,
                 reg614,
                 reg613,
                 reg612,
                 reg611,
                 reg610,
                 reg609,
                 reg608,
                 reg607,
                 forvar606,
                 reg605,
                 reg604,
                 forvar603,
                 reg602,
                 forvar601,
                 reg600,
                 reg599,
                 reg598,
                 forvar597,
                 forvar596,
                 reg595,
                 reg594,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 reg589,
                 forvar588,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 forvar580,
                 reg579,
                 reg578,
                 forvar577,
                 reg576,
                 reg575,
                 reg574,
                 forvar573,
                 forvar572,
                 reg571,
                 wire154,
                 wire156,
                 wire157,
                 wire158,
                 forvar159,
                 reg160,
                 reg161,
                 reg162,
                 reg163,
                 forvar164,
                 reg165,
                 reg166,
                 reg167,
                 reg168,
                 reg169,
                 forvar170,
                 reg171,
                 reg172,
                 reg173,
                 forvar174,
                 reg175,
                 reg176,
                 forvar177,
                 reg178,
                 reg179,
                 reg180,
                 reg181,
                 reg182,
                 reg183,
                 reg184,
                 reg185,
                 forvar186,
                 reg187,
                 reg188,
                 reg189,
                 forvar190,
                 reg191,
                 wire192,
                 wire525,
                 wire527,
                 wire528,
                 wire529,
                 wire530,
                 forvar531,
                 reg532,
                 reg533,
                 reg534,
                 reg535,
                 reg536,
                 reg537,
                 reg538,
                 reg539,
                 reg540,
                 reg541,
                 reg542,
                 reg543,
                 reg544,
                 reg545,
                 reg531,
                 reg546,
                 reg547,
                 reg548,
                 reg549,
                 reg550,
                 reg551,
                 reg552,
                 reg553,
                 reg554,
                 reg555,
                 reg556,
                 reg557,
                 forvar548,
                 reg558,
                 forvar559,
                 reg560,
                 reg561,
                 reg562,
                 reg563,
                 wire564,
                 wire565,
                 wire566,
                 wire567,
                 wire568,
                 wire569,
                 (1'h0)};
  module47 modinst155 (.wire50(wire42), .clk(clk), .wire49(wire44), .wire51(wire43), .y(wire154), .wire48(wire45), .wire52(wire46));
  assign wire156 = $unsigned(wire43);
  assign wire157 = "G";
  assign wire158 = $signed("XbqMnE6XSoRS");
  always
    @(posedge clk) begin
      for (forvar159 = (1'h0); (forvar159 < (3'h4)); forvar159 = (forvar159 + (1'h1)))
        begin
          reg160 <= wire154;
          if (((($unsigned(wire43[(2'h2):(2'h2)]) > wire45[(4'hd):(2'h2)]) ?
                  (!"0qfvZYILpeNDxnvq") : ((!$signed(wire157)) ?
                      wire43[(3'h4):(3'h4)] : wire44)) ?
              ((wire157[(4'he):(4'hd)] >> "mo") ^ $signed("3tv")) : wire158[(2'h2):(2'h2)]))
            begin
              reg161 <= ((~$unsigned($signed(wire46))) <<< ($unsigned(({wire154,
                          reg160} ?
                      $unsigned(wire158) : (wire42 ? (7'h46) : wire42))) ?
                  "9a5KLM4dmzQx97PO8" : ("xuYwEeZEIBkT8" ?
                      ((|wire44) ?
                          wire154[(4'hb):(1'h1)] : $signed(wire42)) : $unsigned((~&wire42)))));
              reg162 <= $unsigned("Ara32i2lS7046uAy9GfOH");
              reg163 <= (wire157[(4'hc):(4'hc)] + (+wire158[(3'h7):(1'h1)]));
            end
          else
            begin
              reg161 <= wire42;
            end
          for (forvar164 = (1'h0); (forvar164 < (2'h2)); forvar164 = (forvar164 + (1'h1)))
            begin
              reg165 <= $signed($unsigned($signed($signed($signed(wire44)))));
              reg166 <= ((^~reg165) ?
                  ($signed((((8'hb3) ? wire156 : wire43) ?
                          (~wire46) : wire42[(4'h8):(4'h8)])) ?
                      wire46[(4'hc):(4'h8)] : reg162[(1'h0):(1'h0)]) : (reg163 > wire44[(3'h7):(3'h4)]));
              reg167 <= "LD";
              reg168 <= $unsigned(((8'h9c) || (((forvar164 ?
                      reg163 : reg163) >> "QDqPnHqhymOpEwH0bRkfJ") ?
                  (!reg166) : "Gk9i")));
              reg169 <= reg161[(4'ha):(1'h1)];
            end
          for (forvar170 = (1'h0); (forvar170 < (1'h1)); forvar170 = (forvar170 + (1'h1)))
            begin
              reg171 = {$signed((!"HxtsNHP6")),
                  $unsigned(((-((7'h48) == wire158)) != (&wire154[(1'h0):(1'h0)])))};
              reg172 <= "kEmFUrN";
              reg173 <= "EVbWBySNh2";
            end
          for (forvar174 = (1'h0); (forvar174 < (2'h2)); forvar174 = (forvar174 + (1'h1)))
            begin
              reg175 <= $signed(reg169);
              reg176 <= wire45[(4'h8):(3'h7)];
            end
        end
      for (forvar177 = (1'h0); (forvar177 < (1'h0)); forvar177 = (forvar177 + (1'h1)))
        begin
          reg178 <= "e0Emt54NW";
          if ((($signed((-(wire156 != reg167))) ?
                  wire157 : reg165[(4'hc):(4'hb)]) ?
              ($signed((8'haf)) ?
                  (($unsigned(forvar174) && $unsigned(reg163)) ?
                      ($signed(wire157) <<< {reg168}) : ($unsigned(reg162) >= "ExSiLy1vTd61")) : (~&(wire46 ?
                      ((8'hb8) >>> reg160) : "DLADxn6PSWJPo"))) : reg168))
            begin
              reg179 <= {reg173[(3'h4):(2'h3)]};
              reg180 <= "Xyu4rEVyNtivg4K";
              reg181 <= forvar177[(4'hd):(2'h3)];
            end
          else
            begin
              reg179 <= (!(8'hbd));
            end
          if ($signed("GbReeK3zf"))
            begin
              reg182 <= (wire154[(1'h0):(1'h0)] ^~ reg168);
            end
          else
            begin
              reg182 <= "ca0";
              reg183 <= "vTFv4DrzyRurgAHo";
              reg184 <= forvar177[(4'hb):(1'h0)];
              reg185 <= $signed($unsigned(forvar177));
            end
          for (forvar186 = (1'h0); (forvar186 < (1'h0)); forvar186 = (forvar186 + (1'h1)))
            begin
              reg187 <= ({$signed($unsigned("YYJfgS3uX5")),
                      ((forvar186 ?
                          wire157[(4'hc):(3'h4)] : {reg172}) >>> $signed((forvar170 ?
                          (7'h45) : wire156)))} ?
                  ((!$unsigned($unsigned(wire44))) << ($signed({(7'h44)}) ?
                      reg180[(2'h2):(2'h2)] : wire156[(3'h6):(3'h5)])) : "");
              reg188 <= reg182;
              reg189 <= {$unsigned($unsigned((-reg175[(5'h14):(4'h8)])))};
            end
          for (forvar190 = (1'h0); (forvar190 < (2'h3)); forvar190 = (forvar190 + (1'h1)))
            begin
              reg191 <= "s";
            end
        end
    end
  assign wire192 = (8'hb3);
  module193 modinst526 (wire525, clk, reg184, wire158, forvar186, reg175);
  assign wire527 = (~($signed(reg162) & forvar177));
  assign wire528 = $signed(reg167);
  assign wire529 = $signed(reg171);
  assign wire530 = reg182[(5'h11):(4'hc)];
  always
    @(posedge clk) begin
      if (((~|reg187) ? $signed("FFCAg24km3K") : reg185))
        begin
          for (forvar531 = (1'h0); (forvar531 < (2'h3)); forvar531 = (forvar531 + (1'h1)))
            begin
              reg532 <= $signed({(~^((|reg189) != reg169[(2'h3):(2'h2)]))});
            end
          if ((~|forvar190[(3'h5):(2'h2)]))
            begin
              reg533 = (~^$unsigned(wire530[(4'hd):(3'h4)]));
              reg534 <= "CsdlWt2bPy";
              reg535 <= reg185[(4'h8):(2'h2)];
              reg536 <= $signed((8'ha9));
            end
          else
            begin
              reg533 <= $unsigned((^$signed($unsigned("yW5DR0GxzJBtN"))));
            end
          if (reg172[(1'h1):(1'h0)])
            begin
              reg537 = ((~&(~^(forvar170 ?
                  ((8'haa) ? (8'hb6) : forvar164) : (reg169 ?
                      reg166 : wire530)))) >= $unsigned("Poed"));
              reg538 <= ($signed("86") | $signed(reg168[(2'h3):(1'h0)]));
            end
          else
            begin
              reg537 <= wire157;
              reg538 <= (~|(~&{reg187}));
              reg539 <= ("" != (reg162[(3'h4):(1'h1)] ?
                  forvar170 : $unsigned((8'ha3))));
              reg540 <= (&reg168[(3'h5):(1'h0)]);
            end
          if (forvar177)
            begin
              reg541 <= (((reg160[(2'h2):(2'h2)] * ("JwDqu5kAgoS03" ~^ (8'hbd))) ?
                  ($unsigned((reg160 >= wire192)) ?
                      $unsigned((reg182 >= reg534)) : $signed((reg532 ?
                          reg183 : wire44))) : ("hUZ9heRY9GM6WkflsCBkN" ?
                      "" : $signed("JorAXBuQ"))) <<< "e5vGx6OiRA6yO1DQCMM7n");
              reg542 <= ("PuSAOoY2O6P" ?
                  $signed((reg535[(4'h9):(1'h0)] ?
                      $signed("K9") : $signed("pmP1oIVcl"))) : "MbuwV5R8ohLliaI7Q8aP");
              reg543 <= {wire46[(4'h9):(3'h6)]};
              reg544 <= ($signed((wire528[(1'h0):(1'h0)] ?
                      $unsigned(wire529) : $signed("696nftZE5y"))) ?
                  reg171[(5'h10):(3'h6)] : (({(wire529 ? wire528 : reg175),
                          reg534} ?
                      forvar186 : $unsigned(wire157)) >>> reg166));
              reg545 <= (^reg171[(4'h9):(1'h1)]);
            end
          else
            begin
              reg541 <= (+"EFk8CUX2Rk6");
              reg542 <= wire158[(3'h5):(2'h2)];
              reg543 <= reg534[(3'h5):(1'h1)];
            end
        end
      else
        begin
          if ((($unsigned({$signed(forvar177)}) ^~ reg178) ?
              {wire528[(1'h1):(1'h1)],
                  $unsigned(((reg543 ? reg161 : (8'hb6)) ?
                      reg182[(4'ha):(4'h8)] : (reg181 ?
                          reg168 : (8'hb3))))} : wire154[(2'h3):(1'h1)]))
            begin
              reg531 <= (^$unsigned($unsigned(forvar164)));
              reg532 <= forvar164[(1'h1):(1'h1)];
              reg533 <= wire529;
              reg534 <= $unsigned("GtrxOzlo5Ue");
              reg535 <= (reg178 - $unsigned(wire46));
            end
          else
            begin
              reg531 <= (forvar170[(2'h3):(2'h2)] > (~&(&$unsigned((forvar531 ?
                  wire525 : (8'ha5))))));
            end
          if (reg161[(1'h1):(1'h0)])
            begin
              reg536 <= $signed($unsigned({"7C8Cvu3t9d"}));
            end
          else
            begin
              reg536 <= reg165[(5'h10):(5'h10)];
            end
          reg537 <= $signed($unsigned(reg160[(3'h4):(1'h0)]));
          reg538 = ("X7yyaS91lfcoeI" ?
              (&"qyukvFu7xdEavTsBuAU") : wire158[(4'ha):(3'h4)]);
        end
      reg546 <= reg185[(1'h1):(1'h1)];
      reg547 <= ($unsigned($unsigned(((~reg188) ?
              $signed(reg532) : ((7'h43) ? forvar177 : reg532)))) ?
          (wire527 * ($signed($signed(wire45)) & forvar174)) : ((~^"LPbhNsymm") ?
              wire154[(3'h6):(3'h5)] : {reg173, reg160[(1'h1):(1'h1)]}));
      if ($unsigned((reg160 <<< "IoN5B")))
        begin
          if ($unsigned(("QXLd7" || reg180[(4'h8):(2'h2)])))
            begin
              reg548 <= forvar159;
              reg549 <= reg183;
              reg550 = wire527[(2'h3):(2'h2)];
              reg551 = $signed(wire156[(3'h5):(1'h1)]);
              reg552 <= $unsigned((~^reg542[(1'h0):(1'h0)]));
            end
          else
            begin
              reg548 <= wire154[(3'h5):(3'h5)];
              reg549 <= $unsigned(reg543);
            end
          if ($signed((((~^$unsigned(wire43)) * wire46) > "343cXy4aIcf")))
            begin
              reg553 <= $unsigned("okl7Z5awvRKNgo1cdV3HcN");
            end
          else
            begin
              reg553 <= "mQM9l";
              reg554 <= $unsigned({($unsigned((reg178 >>> reg178)) == $unsigned("")),
                  (~"DCNfKHQfzusPvalwpBUSV")});
            end
          if ($unsigned(reg191))
            begin
              reg555 <= reg532;
              reg556 = ("PmbSBzABRaCKdZPY4" ?
                  forvar174[(4'h9):(1'h0)] : {reg179[(1'h1):(1'h0)]});
              reg557 <= reg543[(1'h0):(1'h0)];
            end
          else
            begin
              reg555 <= (~&reg540);
              reg556 = (8'h9e);
            end
        end
      else
        begin
          for (forvar548 = (1'h0); (forvar548 < (1'h0)); forvar548 = (forvar548 + (1'h1)))
            begin
              reg549 <= $signed((reg541 < ($signed((forvar159 ?
                      reg557 : (8'hbc))) ?
                  reg167 : $unsigned("nue3dQ8sm01VP2JyYg"))));
              reg550 <= reg191;
              reg551 <= $signed($signed((reg188[(4'ha):(4'h8)] ?
                  {$unsigned(reg544), {wire528, wire525}} : reg166)));
              reg552 <= wire42;
              reg553 <= $unsigned($unsigned(($signed(forvar174) ^~ $signed(forvar164))));
            end
          if (wire192)
            begin
              reg554 <= "ggJOHeu2fYpA08keYu";
              reg555 <= $signed(("3liIvkRkIhk3L7BEHncrUJ" < {(((8'h9e) ?
                      reg533 : reg554) & wire156),
                  $unsigned((~wire527))}));
              reg556 <= ((^("QGgB2JuHROK93w" ?
                      reg555 : "pwibB1UkUo5RkClQBT4C3")) ?
                  "Q" : (("zQFyVID5q" && $signed((~(8'h9d)))) ?
                      $signed({wire154, (^~(8'ha1))}) : "sZLUbIu"));
              reg557 <= "YuytOYRks";
              reg558 <= "GgPV61166C";
            end
          else
            begin
              reg554 = (8'haf);
              reg555 = (|(!reg191[(3'h6):(3'h6)]));
              reg556 <= $signed((^(^~$signed(reg189))));
              reg557 <= wire528;
              reg558 <= ((~&forvar170) != "eLAL");
            end
          for (forvar559 = (1'h0); (forvar559 < (2'h2)); forvar559 = (forvar559 + (1'h1)))
            begin
              reg560 <= $unsigned(("RO" ~^ $signed("lXX2swno3nSR7VWJsv")));
              reg561 <= ((!($signed(reg171[(4'h8):(4'h8)]) ^ "nTnTGUN")) ?
                  (8'hae) : ({reg185} && $unsigned(reg545[(3'h6):(1'h0)])));
              reg562 <= "EavfvvCpK";
              reg563 <= (~&(|(~"MgTBLpKeuirAK")));
            end
        end
    end
  assign wire564 = $unsigned("y7UNKipMSb1pirqTX11");
  assign wire565 = wire46[(3'h5):(3'h4)];
  assign wire566 = (~^reg191);
  assign wire567 = "yLKNH5yv4HUdHB8zgX";
  assign wire568 = $unsigned($unsigned($unsigned(("rC" << reg532))));
  module438 modinst570 (.wire442(reg538), .clk(clk), .y(wire569), .wire440(reg556), .wire443(wire43), .wire439(forvar159), .wire441(forvar190));
  always
    @(posedge clk) begin
      reg571 = $unsigned(reg541[(4'ha):(3'h4)]);
      for (forvar572 = (1'h0); (forvar572 < (1'h0)); forvar572 = (forvar572 + (1'h1)))
        begin
          for (forvar573 = (1'h0); (forvar573 < (1'h1)); forvar573 = (forvar573 + (1'h1)))
            begin
              reg574 = "4G8Y5H1ozK6Mr";
            end
          if (reg179[(2'h2):(1'h1)])
            begin
              reg575 <= "OSEdubwt7mJaSWodXNeFN";
              reg576 <= reg183[(3'h5):(2'h3)];
            end
          else
            begin
              reg575 <= ($signed((!(^~(reg553 >= wire46)))) ?
                  "I1cRr9luYNDt9hbQ" : (~^($signed(reg563[(5'h10):(4'hb)]) ?
                      ((wire564 ?
                          reg171 : reg553) << reg562[(2'h2):(1'h1)]) : (+wire44))));
              reg576 <= ((^{forvar573[(1'h1):(1'h1)]}) ?
                  reg531 : {$signed(((reg541 << reg175) <<< (&reg160)))});
            end
          for (forvar577 = (1'h0); (forvar577 < (2'h3)); forvar577 = (forvar577 + (1'h1)))
            begin
              reg578 <= "ZW";
            end
          reg579 <= {(reg556 ?
                  $signed("cFE3BUXr") : $unsigned("mq96N6XnuxhtKkn3"))};
        end
      for (forvar580 = (1'h0); (forvar580 < (1'h1)); forvar580 = (forvar580 + (1'h1)))
        begin
          if (($signed((({reg571, reg575} & $signed(reg191)) ?
                  "AGUDctn" : reg551[(3'h4):(2'h3)])) ?
              reg540 : $signed(("Bi" >>> ((^reg575) <= "4BW")))))
            begin
              reg581 <= ($unsigned($unsigned(reg172[(2'h2):(1'h0)])) ~^ reg574[(3'h5):(3'h5)]);
              reg582 = reg562[(3'h4):(2'h2)];
            end
          else
            begin
              reg581 <= "4QQ";
              reg582 <= ("9IbEKDgdR3bUADc8yM" << forvar164);
              reg583 <= (((7'h48) >= "D") ?
                  "Jiy1Xs7CgDAe" : (~wire565[(4'hc):(3'h5)]));
            end
          if (($unsigned({{"JeZ99"}}) ?
              ((-reg560[(2'h3):(2'h3)]) > forvar170) : reg173))
            begin
              reg584 <= (^reg546);
            end
          else
            begin
              reg584 <= $signed((((8'hbe) >= reg561) ?
                  $signed($unsigned($signed(reg189))) : ($signed($unsigned(reg165)) ?
                      reg571[(3'h5):(1'h0)] : (|(~|reg532)))));
              reg585 <= "JuN1V9iqp15rd";
              reg586 = "";
              reg587 = (+"LK4hAuDOdBPgJTkCpr");
            end
        end
      for (forvar588 = (1'h0); (forvar588 < (2'h3)); forvar588 = (forvar588 + (1'h1)))
        begin
          reg589 <= reg160;
          if ($unsigned(reg183))
            begin
              reg590 <= (("tJT1PExEvsIdxvsi0fabxu" <= ("WBztq" < "gXGBm4zg")) ^ ($signed(wire528[(1'h1):(1'h0)]) ?
                  (($signed(forvar170) ?
                      (reg180 ^ reg546) : $signed(reg166)) << {$signed(wire157),
                      $signed(reg583)}) : (reg166[(3'h4):(1'h0)] || ($signed(wire528) ?
                      $signed(reg561) : (~reg166)))));
              reg591 <= (reg175 ? $signed((~&"wMg")) : reg539[(1'h0):(1'h0)]);
              reg592 <= $signed("n8f9VMO1");
              reg593 <= (&forvar159[(2'h3):(1'h1)]);
            end
          else
            begin
              reg590 <= (reg183 ? reg571 : (reg545 <= (~&$unsigned(reg162))));
              reg591 <= (!reg160[(2'h2):(1'h1)]);
              reg592 <= (8'hb8);
              reg593 <= reg185;
            end
          reg594 <= (($unsigned($signed(wire564[(4'hd):(3'h6)])) ^ ((~^(reg178 ?
                  reg579 : reg552)) ?
              ($unsigned(reg173) ?
                  (~&reg590) : $unsigned(forvar186)) : {(reg571 ?
                      reg548 : reg179)})) | $unsigned((($signed(reg183) < (reg187 ?
              (8'h9e) : wire192)) - (8'h9f))));
          reg595 <= reg166;
        end
      for (forvar596 = (1'h0); (forvar596 < (2'h3)); forvar596 = (forvar596 + (1'h1)))
        begin
          for (forvar597 = (1'h0); (forvar597 < (1'h0)); forvar597 = (forvar597 + (1'h1)))
            begin
              reg598 <= $unsigned(({(~$unsigned(reg575))} ^ "fGXX9Tyl9m6zUBhSa"));
            end
          reg599 = "K5XQaZ";
        end
    end
  always
    @(posedge clk) begin
      reg600 <= "SC6gN7klbZ";
      for (forvar601 = (1'h0); (forvar601 < (2'h2)); forvar601 = (forvar601 + (1'h1)))
        begin
          reg602 <= wire530[(4'h8):(4'h8)];
          for (forvar603 = (1'h0); (forvar603 < (2'h3)); forvar603 = (forvar603 + (1'h1)))
            begin
              reg604 <= $signed(forvar597[(1'h0):(1'h0)]);
              reg605 <= $signed("Nu6Eknhz7");
            end
          for (forvar606 = (1'h0); (forvar606 < (2'h3)); forvar606 = (forvar606 + (1'h1)))
            begin
              reg607 <= (reg556[(4'h8):(4'h8)] ^ (~^reg589));
              reg608 <= reg595[(4'he):(3'h7)];
            end
          if (("isGyBWr15ItA" >= (("WT2xMZI44k3n" > ($unsigned(reg576) ?
                  (+(8'hb8)) : "kNS07dtEeFp")) ?
              forvar548[(4'hd):(1'h1)] : wire530)))
            begin
              reg609 <= "eyBRKT";
            end
          else
            begin
              reg609 = (!$signed(""));
              reg610 <= forvar606[(2'h3):(2'h3)];
              reg611 <= reg609[(4'ha):(4'h8)];
              reg612 = $unsigned((((reg535[(4'h9):(3'h7)] ?
                  $unsigned(reg561) : "AyIql5gY93EyGmMESzW") ^ (((8'hb1) == reg188) ?
                  (reg594 <<< (8'hb7)) : (reg183 != reg181))) ^~ reg178[(1'h0):(1'h0)]));
              reg613 <= $unsigned((&$signed({{reg179}})));
            end
          reg614 = {"2Ma3Oz4ENSDeFMza8vitXW"};
        end
      for (forvar615 = (1'h0); (forvar615 < (2'h2)); forvar615 = (forvar615 + (1'h1)))
        begin
          reg616 <= $unsigned($signed($signed({reg614[(5'h11):(1'h0)],
              ((8'hae) - forvar190)})));
          reg617 <= $unsigned($signed((reg602 ? "KTe0L" : "6188CUKO4LGYB")));
        end
    end
  assign wire618 = "mD6CGuvTWweYD1KoInAkR";
  always
    @(posedge clk) begin
      reg619 <= ((~&{({forvar580, forvar601} ?
              (reg556 ? reg599 : (8'hae)) : (reg552 ?
                  reg591 : reg585))}) | ((reg541[(1'h1):(1'h0)] ?
          forvar597[(5'h11):(1'h0)] : {$signed(reg585)}) == (($unsigned(reg563) ?
          (8'hb3) : (reg592 == reg168)) << $signed((^~wire154)))));
      if ($signed("wbHXdV8ZT"))
        begin
          for (forvar620 = (1'h0); (forvar620 < (2'h2)); forvar620 = (forvar620 + (1'h1)))
            begin
              reg621 <= {reg604[(3'h5):(2'h2)],
                  (((forvar573 ?
                          reg554 : (forvar573 ?
                              reg544 : reg554)) < forvar615[(2'h2):(2'h2)]) ?
                      ({((8'hbf) ?
                              forvar186 : forvar572)} >>> ((~|forvar596) & (7'h45))) : reg612[(2'h3):(2'h3)])};
              reg622 <= {"EgioR", "q2m73Buri3F5Th8lGF"};
              reg623 <= "oPIe0OgOYPxF6pe";
              reg624 <= "OATubDsUUu6KEYm0w";
              reg625 <= (^~$signed(forvar588[(3'h5):(1'h1)]));
            end
          if (((~^reg604) ?
              "Mbp6u0xhLJGeTuNUk7M" : $signed($signed((~&{reg594, reg547})))))
            begin
              reg626 <= (($unsigned(((|(8'hb6)) ?
                      (reg561 | reg556) : $signed(wire530))) ?
                  ((reg535[(2'h2):(1'h1)] ?
                          reg536 : (wire567 ? wire45 : reg179)) ?
                      wire192[(1'h1):(1'h0)] : $unsigned({reg531})) : $signed(reg616[(1'h1):(1'h1)])) * $signed(wire569));
              reg627 = "rbKx2DclBZh";
              reg628 <= $signed("y");
              reg629 <= $signed((~($unsigned((reg160 ?
                  reg552 : reg185)) ^ (^(!reg556)))));
              reg630 = ("r" << $signed(forvar190[(4'h8):(3'h4)]));
            end
          else
            begin
              reg626 <= {"",
                  ((&reg191[(3'h5):(2'h2)]) >>> "OmmZuAFUChlATiA4w3")};
              reg627 <= (reg574[(1'h1):(1'h0)] & reg592[(4'h9):(2'h2)]);
              reg628 <= $signed({wire44[(2'h3):(2'h2)]});
              reg629 <= {reg183[(3'h7):(3'h4)],
                  ("IR6IW" ?
                      "zvm5y7O0HhEAoD7aHEZ" : ($signed((reg609 ~^ forvar606)) && "R"))};
              reg630 <= ($unsigned((("cplTOXtoY" ?
                      (reg185 ?
                          reg583 : reg551) : "B2WX4gSKeVL8X") < (+{forvar596,
                      (8'hbf)}))) ?
                  $unsigned(wire618[(2'h2):(1'h0)]) : reg160[(2'h2):(2'h2)]);
            end
          reg631 <= forvar573;
          reg632 <= (($unsigned(($signed(reg160) ?
                  reg594[(3'h4):(1'h0)] : forvar596[(4'h9):(1'h0)])) ?
              $signed({(8'ha5)}) : $unsigned(((reg191 ? reg593 : reg191) ?
                  "tnaZ" : "RZNgTWH"))) << reg583);
        end
      else
        begin
          for (forvar620 = (1'h0); (forvar620 < (2'h3)); forvar620 = (forvar620 + (1'h1)))
            begin
              reg621 <= ($unsigned((($signed(reg625) ?
                          (reg163 | forvar559) : "9g27g8GFiQ") ?
                      "VVIAI" : reg188[(1'h1):(1'h0)])) ?
                  (($signed((wire46 >= forvar615)) | reg612[(1'h0):(1'h0)]) ?
                      ($signed({reg561,
                          reg571}) * "pxCK46GfsUZ0L1Hx") : $signed($unsigned("UDyDGIIKUMi"))) : (~reg551));
              reg622 <= {{reg533, reg183}};
              reg623 <= "azrT";
            end
          reg624 <= reg538[(4'h9):(4'h9)];
          for (forvar625 = (1'h0); (forvar625 < (1'h1)); forvar625 = (forvar625 + (1'h1)))
            begin
              reg626 <= $signed((((8'ha9) <= ($unsigned(wire564) ?
                      (^reg181) : (wire530 ? wire158 : forvar164))) ?
                  (+"zGsIOxblzD") : reg534[(3'h7):(1'h0)]));
              reg627 <= "P3CZprQszi";
              reg628 = $signed("glMZs3vhsDOeGa");
            end
        end
      reg633 <= wire530;
      for (forvar634 = (1'h0); (forvar634 < (1'h0)); forvar634 = (forvar634 + (1'h1)))
        begin
          reg635 <= "";
          if ((^~$unsigned($unsigned($signed((8'haf))))))
            begin
              reg636 <= (($unsigned(reg549) << ({forvar596} ?
                      reg578 : ("xesfB" ?
                          $signed(forvar577) : $unsigned(reg182)))) ?
                  (wire527 * reg584) : {(~|(wire525 >>> reg180[(4'he):(4'h8)]))});
              reg637 <= reg176;
              reg638 <= (-"C2Dc1mZKYl");
            end
          else
            begin
              reg636 <= {$signed(($unsigned(reg582) ^~ ((forvar615 ?
                      (8'h9f) : (8'h9f)) <= reg173)))};
              reg637 <= (^~reg539[(5'h17):(3'h7)]);
              reg638 <= $signed(wire567[(5'h13):(4'he)]);
              reg639 <= reg532[(2'h2):(2'h2)];
              reg640 <= reg537;
            end
          for (forvar641 = (1'h0); (forvar641 < (1'h1)); forvar641 = (forvar641 + (1'h1)))
            begin
              reg642 <= "";
              reg643 <= wire157[(1'h0):(1'h0)];
              reg644 <= $unsigned((8'ha1));
              reg645 <= "t9INNU1YOsR7MywkCES";
            end
        end
      if ((~(^~$unsigned(wire158))))
        begin
          reg646 <= ("zSMPtk2fcNQFASxKslwei" + reg180);
          if ($unsigned((reg547 ?
              reg543[(2'h2):(2'h2)] : (!{reg180[(1'h0):(1'h0)],
                  ((7'h42) ? (7'h40) : reg630)}))))
            begin
              reg647 <= {"NxtycVXu", $signed($signed($signed(reg547)))};
              reg648 <= (~^(~wire43));
              reg649 <= $unsigned((~|(reg630[(4'hd):(3'h6)] ?
                  reg562 : $unsigned((reg540 * forvar177)))));
            end
          else
            begin
              reg647 <= (reg625 ?
                  ((|reg602) - ($unsigned(reg587) ?
                      (((8'hb8) ? reg182 : reg640) ?
                          $unsigned(reg552) : (reg542 ?
                              forvar577 : wire564)) : reg553)) : ($unsigned(($unsigned(reg167) != $unsigned(reg647))) & $signed($signed($unsigned(wire565)))));
              reg648 <= "MtOFxCnP4OE3MWSADF440";
            end
          for (forvar650 = (1'h0); (forvar650 < (2'h2)); forvar650 = (forvar650 + (1'h1)))
            begin
              reg651 <= ("u5sHwt9rTyKc" >>> ((&wire154[(4'hf):(2'h2)]) ?
                  (^~((+reg649) ?
                      $unsigned(reg553) : (^~(8'ha2)))) : $signed(reg604[(2'h2):(2'h2)])));
            end
          for (forvar652 = (1'h0); (forvar652 < (1'h1)); forvar652 = (forvar652 + (1'h1)))
            begin
              reg653 <= (~|$unsigned($unsigned(reg576)));
              reg654 <= (~&{$unsigned($unsigned((|reg647))),
                  {reg605,
                      ((reg167 ^~ wire569) ?
                          $signed(reg623) : reg538[(4'hb):(4'h9)])}});
              reg655 <= "AQMXLFVqmNsBPzA1vvw";
              reg656 <= reg629;
              reg657 <= $signed((forvar573 ? reg595 : wire569));
            end
        end
      else
        begin
          for (forvar646 = (1'h0); (forvar646 < (2'h3)); forvar646 = (forvar646 + (1'h1)))
            begin
              reg647 <= $signed(($signed((forvar625[(4'ha):(4'ha)] + (reg611 != reg533))) ?
                  (&reg608[(1'h1):(1'h1)]) : "zT6ackPQXWS1oLny1hUFH"));
              reg648 <= reg591[(2'h3):(2'h3)];
              reg649 <= "AMRrSAeEnfOfoA3D";
            end
          reg650 <= forvar531[(1'h0):(1'h0)];
          for (forvar651 = (1'h0); (forvar651 < (1'h0)); forvar651 = (forvar651 + (1'h1)))
            begin
              reg652 = $signed(reg575[(3'h7):(3'h7)]);
              reg653 <= reg175;
              reg654 <= (~^$signed((forvar559 ?
                  $signed(reg537) : $signed(reg166[(3'h7):(1'h0)]))));
              reg655 <= (forvar577 != reg163[(5'h13):(4'hc)]);
              reg656 <= reg581[(2'h2):(2'h2)];
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module193  (y, clk, wire194, wire195, wire196, wire197);
  output wire [(32'h657):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire194;
  input wire [(4'hb):(1'h0)] wire195;
  input wire [(2'h2):(1'h0)] wire196;
  input wire signed [(5'h13):(1'h0)] wire197;
  reg signed [(4'h8):(1'h0)] reg524 = (1'h0);
  reg [(4'h8):(1'h0)] reg523 = (1'h0);
  reg [(4'he):(1'h0)] reg522 = (1'h0);
  reg [(4'hd):(1'h0)] reg521 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg520 = (1'h0);
  wire [(5'h11):(1'h0)] wire391;
  wire [(5'h14):(1'h0)] wire351;
  wire signed [(5'h14):(1'h0)] wire349;
  reg signed [(3'h4):(1'h0)] reg312 = (1'h0);
  reg [(4'hb):(1'h0)] reg311 = (1'h0);
  reg [(4'hd):(1'h0)] reg307 = (1'h0);
  reg [(2'h2):(1'h0)] reg310 = (1'h0);
  reg [(2'h2):(1'h0)] reg309 = (1'h0);
  reg [(4'hc):(1'h0)] reg308 = (1'h0);
  reg [(4'he):(1'h0)] forvar307 = (1'h0);
  reg [(5'h13):(1'h0)] reg306 = (1'h0);
  reg [(4'hd):(1'h0)] reg305 = (1'h0);
  reg [(5'h10):(1'h0)] reg290 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg304 = (1'h0);
  reg [(4'hc):(1'h0)] reg303 = (1'h0);
  reg [(2'h3):(1'h0)] reg302 = (1'h0);
  reg [(4'hc):(1'h0)] reg301 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg300 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg299 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg298 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg297 = (1'h0);
  reg [(5'h11):(1'h0)] reg296 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg295 = (1'h0);
  reg [(4'hf):(1'h0)] reg294 = (1'h0);
  reg [(5'h14):(1'h0)] forvar293 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg292 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg291 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar290 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar287 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg283 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg278 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg289 = (1'h0);
  reg [(4'ha):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg287 = (1'h0);
  reg [(3'h7):(1'h0)] reg286 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg285 = (1'h0);
  reg [(2'h3):(1'h0)] reg284 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar283 = (1'h0);
  reg [(5'h10):(1'h0)] reg282 = (1'h0);
  reg [(4'h8):(1'h0)] reg281 = (1'h0);
  reg [(4'h9):(1'h0)] reg280 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg279 = (1'h0);
  reg [(3'h5):(1'h0)] forvar278 = (1'h0);
  reg signed [(4'he):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg276 = (1'h0);
  reg [(3'h6):(1'h0)] reg275 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar274 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire273;
  wire signed [(2'h3):(1'h0)] wire272;
  wire signed [(5'h12):(1'h0)] wire271;
  reg [(4'hb):(1'h0)] reg270 = (1'h0);
  reg [(5'h11):(1'h0)] reg269 = (1'h0);
  reg [(5'h15):(1'h0)] reg268 = (1'h0);
  reg [(3'h6):(1'h0)] reg267 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar266 = (1'h0);
  reg [(2'h3):(1'h0)] reg265 = (1'h0);
  reg [(4'hb):(1'h0)] reg264 = (1'h0);
  reg [(4'hb):(1'h0)] forvar263 = (1'h0);
  reg [(5'h10):(1'h0)] reg262 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg261 = (1'h0);
  reg [(5'h11):(1'h0)] reg260 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg259 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg258 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg253 = (1'h0);
  reg [(5'h16):(1'h0)] reg257 = (1'h0);
  reg [(4'hd):(1'h0)] reg256 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg255 = (1'h0);
  reg [(5'h13):(1'h0)] reg254 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar253 = (1'h0);
  reg [(2'h2):(1'h0)] reg252 = (1'h0);
  wire [(4'hd):(1'h0)] wire251;
  wire [(4'hb):(1'h0)] wire198;
  wire signed [(5'h11):(1'h0)] wire199;
  wire signed [(3'h6):(1'h0)] wire249;
  wire [(5'h14):(1'h0)] wire393;
  reg signed [(3'h4):(1'h0)] reg394 = (1'h0);
  reg [(5'h16):(1'h0)] forvar395 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg396 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg397 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar398 = (1'h0);
  reg [(5'h11):(1'h0)] reg399 = (1'h0);
  reg [(2'h3):(1'h0)] reg400 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg401 = (1'h0);
  reg [(4'hd):(1'h0)] reg402 = (1'h0);
  reg [(3'h7):(1'h0)] reg403 = (1'h0);
  reg signed [(4'he):(1'h0)] reg404 = (1'h0);
  reg [(3'h5):(1'h0)] reg405 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg406 = (1'h0);
  reg [(4'he):(1'h0)] reg407 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg408 = (1'h0);
  reg [(4'hc):(1'h0)] reg409 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg410 = (1'h0);
  reg [(4'he):(1'h0)] reg411 = (1'h0);
  reg [(3'h7):(1'h0)] forvar400 = (1'h0);
  reg [(4'hf):(1'h0)] forvar412 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg413 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg414 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg415 = (1'h0);
  reg [(4'hd):(1'h0)] reg416 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg417 = (1'h0);
  reg [(3'h7):(1'h0)] reg418 = (1'h0);
  reg [(3'h7):(1'h0)] reg419 = (1'h0);
  reg [(2'h2):(1'h0)] reg420 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg421 = (1'h0);
  reg [(5'h13):(1'h0)] forvar422 = (1'h0);
  reg [(5'h10):(1'h0)] reg423 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg424 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg425 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg426 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg427 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar428 = (1'h0);
  reg [(5'h10):(1'h0)] reg429 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg430 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar431 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg432 = (1'h0);
  reg [(3'h7):(1'h0)] reg433 = (1'h0);
  reg [(5'h13):(1'h0)] reg434 = (1'h0);
  reg [(5'h10):(1'h0)] reg435 = (1'h0);
  wire signed [(4'he):(1'h0)] wire436;
  wire signed [(2'h2):(1'h0)] wire437;
  wire signed [(4'h8):(1'h0)] wire518;
  assign y = {reg524,
                 reg523,
                 reg522,
                 reg521,
                 reg520,
                 wire391,
                 wire351,
                 wire349,
                 reg312,
                 reg311,
                 reg307,
                 reg310,
                 reg309,
                 reg308,
                 forvar307,
                 reg306,
                 reg305,
                 reg290,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 reg298,
                 reg297,
                 reg296,
                 reg295,
                 reg294,
                 forvar293,
                 reg292,
                 reg291,
                 forvar290,
                 forvar287,
                 reg283,
                 reg278,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 forvar283,
                 reg282,
                 reg281,
                 reg280,
                 reg279,
                 forvar278,
                 reg277,
                 reg276,
                 reg275,
                 forvar274,
                 wire273,
                 wire272,
                 wire271,
                 reg270,
                 reg269,
                 reg268,
                 reg267,
                 forvar266,
                 reg265,
                 reg264,
                 forvar263,
                 reg262,
                 reg261,
                 reg260,
                 reg259,
                 reg258,
                 reg253,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 forvar253,
                 reg252,
                 wire251,
                 wire198,
                 wire199,
                 wire249,
                 wire393,
                 reg394,
                 forvar395,
                 reg396,
                 reg397,
                 forvar398,
                 reg399,
                 reg400,
                 reg401,
                 reg402,
                 reg403,
                 reg404,
                 reg405,
                 reg406,
                 reg407,
                 reg408,
                 reg409,
                 reg410,
                 reg411,
                 forvar400,
                 forvar412,
                 reg413,
                 reg414,
                 reg415,
                 reg416,
                 reg417,
                 reg418,
                 reg419,
                 reg420,
                 reg421,
                 forvar422,
                 reg423,
                 reg424,
                 reg425,
                 reg426,
                 reg427,
                 forvar428,
                 reg429,
                 reg430,
                 forvar431,
                 reg432,
                 reg433,
                 reg434,
                 reg435,
                 wire436,
                 wire437,
                 wire518,
                 (1'h0)};
  assign wire198 = (wire194[(2'h3):(2'h2)] ^~ ($signed($signed("koB5MfJFpQ")) ?
                       (+$unsigned((~^(8'hab)))) : ""));
  assign wire199 = {(wire198[(1'h0):(1'h0)] ?
                           $signed((8'hb8)) : ((!wire198) * wire194))};
  module200 modinst250 (wire249, clk, wire195, wire199, wire197, wire194, wire198);
  assign wire251 = $unsigned(($unsigned($signed(wire249[(2'h3):(2'h3)])) <<< ((wire196[(1'h1):(1'h1)] ^ (8'hbb)) ?
                       wire197[(4'hb):(4'h9)] : wire198[(1'h1):(1'h0)])));
  always
    @(posedge clk) begin
      if (($signed(((|wire249) ?
              (&(wire194 + wire194)) : $unsigned({wire197, wire197}))) ?
          {wire197} : wire198[(1'h0):(1'h0)]))
        begin
          reg252 <= (^~(&$signed((8'hb9))));
          for (forvar253 = (1'h0); (forvar253 < (2'h3)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 <= "qNafMyrTJ";
              reg255 <= ("R4NLIg" < "z");
              reg256 <= $signed("wo0cT5Sfwdnqk");
            end
          reg257 = $signed(reg252);
        end
      else
        begin
          if (("zG8bO7T1fohZTtx0R1Z" ^ $signed(wire249)))
            begin
              reg252 <= ((&{((~&wire194) ?
                      wire199 : wire199)}) ^ ({$signed((wire194 ?
                      reg252 : wire249)),
                  (reg254[(4'hb):(1'h0)] ?
                      wire199 : wire197[(5'h11):(5'h11)])} - wire195));
            end
          else
            begin
              reg252 <= wire197[(4'hf):(4'he)];
              reg253 <= $unsigned("MI3R1KF7");
              reg254 = reg256[(4'h8):(3'h6)];
            end
          if (($unsigned(((reg256[(4'ha):(4'h9)] ?
                  $unsigned(reg252) : forvar253) && ($unsigned(wire195) < forvar253[(3'h7):(3'h4)]))) ?
              ({(wire251[(1'h1):(1'h1)] ?
                          $signed(wire198) : $unsigned(wire194))} ?
                  (~|$signed((wire196 ?
                      reg253 : wire199))) : {$unsigned((reg252 ?
                          (8'h9e) : wire197))}) : {{reg252[(1'h1):(1'h0)],
                      (reg252[(1'h0):(1'h0)] <= reg257[(5'h16):(3'h5)])}}))
            begin
              reg255 <= ((-($unsigned(wire195) ?
                      ((wire195 << wire195) != wire199) : wire249)) ?
                  {({{wire251}, $signed(reg253)} ?
                          "" : (reg257 ? {reg257} : (~^reg253))),
                      wire195} : $signed(("yD0bJl" >>> "n0Mgf4MV")));
              reg256 <= $signed({$signed($signed({wire251, reg253})),
                  ("8HzaeusX" ?
                      (^~(&wire199)) : (forvar253[(1'h1):(1'h1)] <<< wire249[(1'h0):(1'h0)]))});
            end
          else
            begin
              reg255 <= reg254;
              reg256 <= $unsigned(((8'ha4) ?
                  ("ZVUMfA53DC" ?
                      $signed(((8'ha2) ?
                          wire199 : reg254)) : $signed((-wire196))) : "fm1MSFM5hXSZVyZWq"));
              reg257 = wire196;
              reg258 <= $unsigned((~$unsigned("zbCDO")));
              reg259 <= wire196[(1'h1):(1'h0)];
            end
          if ($signed((!($signed("fdygzOi9IP9LCT4qm7eZs") ?
              $signed($signed(reg257)) : ((7'h40) ? {wire249} : (|reg258))))))
            begin
              reg260 = {(($unsigned("xE0ohlmwvwGYoEvmY5BV") ?
                          ((7'h48) << $unsigned(wire199)) : ($unsigned(wire199) == forvar253[(5'h11):(3'h7)])) ?
                      wire197[(5'h10):(4'hb)] : {({reg259} ?
                              reg257 : $unsigned(reg252)),
                          reg256[(1'h1):(1'h1)]}),
                  {($signed($signed(wire197)) <<< (wire194 >> ((8'ha5) ?
                          reg255 : wire194)))}};
              reg261 <= $signed(((~|(~^(wire195 ?
                  wire196 : (8'ha1)))) && {(reg260[(4'hf):(4'h8)] ?
                      $unsigned(reg260) : reg252)}));
              reg262 = (+$unsigned(wire251));
            end
          else
            begin
              reg260 <= (-{$signed($signed((8'h9c))), "EDBzta7a"});
              reg261 <= reg258;
            end
          for (forvar263 = (1'h0); (forvar263 < (2'h2)); forvar263 = (forvar263 + (1'h1)))
            begin
              reg264 <= ($signed(wire194[(3'h7):(3'h5)]) ?
                  $signed($signed($signed(reg256[(4'h9):(2'h2)]))) : "J0hq6fEQX");
              reg265 <= $signed((wire199 != "E7er8mHt1N9CTc"));
            end
          for (forvar266 = (1'h0); (forvar266 < (2'h3)); forvar266 = (forvar266 + (1'h1)))
            begin
              reg267 <= reg252[(2'h2):(2'h2)];
              reg268 <= $unsigned(forvar266[(2'h3):(2'h2)]);
              reg269 <= ({$unsigned(wire198[(2'h3):(1'h1)]),
                  "mO3kvxrGVqBOfYp"} > {{(^{reg268}),
                      (((8'h9d) ^ forvar253) ?
                          forvar263 : (reg265 && wire195))},
                  ("Z6pMGTeJBkhz4fPLKStwR" > reg253)});
              reg270 = (reg261[(2'h2):(1'h1)] <= reg253[(2'h2):(1'h1)]);
            end
        end
    end
  assign wire271 = (wire195 ?
                       (wire195 ?
                           $unsigned(($unsigned((8'hb6)) ?
                               wire251[(1'h1):(1'h1)] : ((8'ha3) ?
                                   reg257 : reg269))) : (wire194[(1'h0):(1'h0)] ?
                               (^~$signed(wire251)) : reg267)) : reg270);
  assign wire272 = "f0CN4l6HMQ1PFT9gVywr";
  assign wire273 = "p6GXd";
  always
    @(posedge clk) begin
      if ((|"u"))
        begin
          for (forvar274 = (1'h0); (forvar274 < (2'h2)); forvar274 = (forvar274 + (1'h1)))
            begin
              reg275 <= $unsigned(reg254);
              reg276 <= reg275;
              reg277 <= ({"TyfOZo7xm5oMYDEtzo",
                  $unsigned(((wire197 ? reg262 : reg255) ?
                      (reg276 ?
                          reg270 : reg276) : "c9nwt9heTWn"))} >> ({reg260} ?
                  $unsigned($signed((^~wire196))) : (8'hb1)));
            end
          for (forvar278 = (1'h0); (forvar278 < (2'h3)); forvar278 = (forvar278 + (1'h1)))
            begin
              reg279 <= ("CI2Mhqs32UHC" < (($unsigned(wire249[(3'h5):(2'h3)]) >= ((reg261 ^~ reg270) ?
                      wire195[(1'h0):(1'h0)] : reg275)) ?
                  (^(reg260 ?
                      (reg253 + wire194) : "tKyyl7g5Lz3UH9aQre76")) : reg267[(2'h3):(2'h3)]));
              reg280 <= $unsigned("v0lQ5IqbgPEZJmtFnXXSU0");
              reg281 <= "BuD5A";
              reg282 <= ("" ? (|reg268[(5'h13):(4'hf)]) : "e");
            end
          for (forvar283 = (1'h0); (forvar283 < (1'h1)); forvar283 = (forvar283 + (1'h1)))
            begin
              reg284 <= ((reg256[(4'h8):(3'h6)] ? "qkmAOlfhZ" : reg275) ?
                  ((reg269[(4'h9):(3'h5)] >= wire273) ~^ wire194) : ((forvar274[(2'h2):(2'h2)] < forvar263) ?
                      forvar253 : "Azgq"));
            end
          if (wire196[(1'h0):(1'h0)])
            begin
              reg285 = reg252;
            end
          else
            begin
              reg285 <= (~|$signed($signed($signed(reg275[(1'h1):(1'h0)]))));
              reg286 <= $unsigned(reg259);
              reg287 <= (^($unsigned($signed(reg277[(4'h8):(1'h1)])) ?
                  $unsigned(({reg269} && reg254)) : "P3HLtdEC"));
              reg288 = reg261[(3'h4):(1'h1)];
              reg289 <= "3JaIetsSPW";
            end
        end
      else
        begin
          for (forvar274 = (1'h0); (forvar274 < (1'h1)); forvar274 = (forvar274 + (1'h1)))
            begin
              reg275 <= "g8";
              reg276 = ($signed($signed(forvar274)) == reg285[(2'h2):(1'h1)]);
              reg277 <= wire198;
              reg278 <= (reg268[(5'h13):(4'h8)] ~^ (&$signed(reg255[(3'h6):(1'h1)])));
            end
          if ((8'ha6))
            begin
              reg279 <= wire198[(4'h9):(3'h7)];
              reg280 = reg276;
              reg281 <= (8'hb0);
            end
          else
            begin
              reg279 = {(|reg262[(1'h0):(1'h0)])};
              reg280 <= reg256;
            end
          if ((-$signed(reg264)))
            begin
              reg282 <= ({reg253, (~&$signed("PHnoexS0aUlV7tqQ"))} ?
                  $signed($unsigned("cSQspWtO1qEHf8")) : wire194);
              reg283 <= (reg259[(1'h0):(1'h0)] >>> $unsigned((^wire195)));
              reg284 <= $unsigned({(({reg258, forvar283} ?
                      reg281[(2'h2):(1'h1)] : $unsigned((8'hbb))) != ($signed(reg262) ?
                      $unsigned(reg276) : (wire249 ? wire195 : reg253)))});
              reg285 <= wire195[(4'hb):(3'h4)];
            end
          else
            begin
              reg282 <= reg255;
              reg283 <= $signed(reg259);
              reg284 <= $unsigned("d0Gg8VYpxoYGlVC");
              reg285 <= $signed((~|$unsigned((|(+reg258)))));
              reg286 <= ((&$unsigned("LAvhrIllkvvYUMViviX")) ^~ (reg286[(2'h3):(2'h2)] >> ({{reg268,
                      wire271},
                  (&wire197)} == wire199)));
            end
          for (forvar287 = (1'h0); (forvar287 < (3'h4)); forvar287 = (forvar287 + (1'h1)))
            begin
              reg288 <= reg281;
              reg289 <= reg276;
            end
        end
      if (reg257)
        begin
          for (forvar290 = (1'h0); (forvar290 < (1'h1)); forvar290 = (forvar290 + (1'h1)))
            begin
              reg291 <= "4AkxnAnIQx8E6MSUVfh";
              reg292 = {"2I4llACo8wbvH4ydTXERa"};
            end
          for (forvar293 = (1'h0); (forvar293 < (3'h4)); forvar293 = (forvar293 + (1'h1)))
            begin
              reg294 <= "EurpGoBMLWKCuPo";
              reg295 <= forvar293[(3'h5):(1'h0)];
              reg296 <= forvar283[(4'hf):(2'h2)];
              reg297 = ($signed($unsigned($signed($signed((8'hb7))))) ?
                  {wire194[(5'h12):(3'h5)],
                      (((reg259 - wire271) ?
                          wire197 : (&reg265)) >>> $unsigned($signed(forvar293)))} : (~|({(^~wire249)} << (((8'hb2) > wire194) ?
                      $signed(wire197) : wire199))));
            end
          if ((-$signed($signed((^~$unsigned(reg295))))))
            begin
              reg298 <= $unsigned((($signed(reg286[(2'h2):(1'h1)]) & $signed(forvar263)) ?
                  reg291[(1'h1):(1'h0)] : {$unsigned($signed(forvar287))}));
              reg299 <= (^~(8'hbe));
              reg300 <= reg289;
              reg301 <= reg283;
              reg302 <= $unsigned($signed({("Db6" - (~reg279))}));
            end
          else
            begin
              reg298 <= {"Q"};
              reg299 <= "JdrY7KCNqtENZ7";
              reg300 <= $signed({""});
            end
          reg303 <= "teqw";
          reg304 <= "kl7EeBIvzt3m27Xb";
        end
      else
        begin
          reg290 <= $signed(($unsigned($signed(((8'hb1) ?
                  forvar278 : wire194))) ?
              ($signed(reg252[(1'h0):(1'h0)]) < "") : reg259));
        end
      if ((&forvar263))
        begin
          if ($signed("AbGbpaVa5xewqx"))
            begin
              reg305 <= reg285[(4'ha):(4'h8)];
              reg306 = (forvar290 <= {($unsigned("H8ge0") ?
                      reg297 : $unsigned((-reg267))),
                  ({wire249[(2'h2):(1'h0)],
                      "892T3WnbLBhfEsH"} > (~(reg262 << (8'h9c))))});
            end
          else
            begin
              reg305 = (~$unsigned((|forvar263[(1'h1):(1'h0)])));
            end
          for (forvar307 = (1'h0); (forvar307 < (2'h3)); forvar307 = (forvar307 + (1'h1)))
            begin
              reg308 <= "blqO86pQBNo";
              reg309 <= forvar283[(3'h7):(1'h0)];
            end
          reg310 <= $signed($signed((forvar287 <= ((&reg256) > (reg275 >>> reg283)))));
        end
      else
        begin
          if (reg295[(4'hf):(4'ha)])
            begin
              reg305 <= reg295[(5'h10):(3'h7)];
            end
          else
            begin
              reg305 <= {wire272, {"NPt", forvar278[(1'h0):(1'h0)]}};
              reg306 <= $unsigned($signed(wire273));
              reg307 = (~"Ogukb6192H3PJb");
            end
          if ({(|reg258),
              ((~|(reg300[(4'he):(3'h6)] ^ (reg262 ? reg299 : forvar307))) ?
                  reg270[(1'h0):(1'h0)] : "ziwbQZgEVeVT")})
            begin
              reg308 <= (7'h48);
              reg309 <= {(|"TK17Ur3whfU0pnwU"), reg307[(3'h4):(1'h0)]};
              reg310 <= (("TNszAcXezTbmVFq2ko" ?
                      (((wire271 ? reg306 : (7'h44)) < (reg289 ?
                          wire196 : wire273)) ^~ "WYrlMkhSMqN76J") : ("Ww9w01Y36gywwqZWB6cq" - $signed({wire249}))) ?
                  (~|(($unsigned((7'h47)) >= (reg298 ~^ reg308)) ?
                      (7'h44) : $signed({forvar253,
                          reg281}))) : ($signed(((reg276 || wire251) ?
                          {reg296} : ((8'ha7) != reg295))) ?
                      "cbGs9Xbhsy5Tvt50F72TqI" : ("OY2chbvU8T6CzW" ?
                          $signed("zWaw7awNPLHyx9") : reg270[(3'h6):(3'h6)])));
              reg311 <= reg259[(2'h3):(1'h1)];
              reg312 <= ($unsigned(((8'hba) ?
                      ("IkkiYkiz" - $unsigned(wire195)) : (reg282[(3'h6):(1'h1)] ?
                          (wire195 != reg290) : (&reg261)))) ?
                  $unsigned($unsigned((8'hb6))) : $signed("1iO2gtUWmNtAtacqB4"));
            end
          else
            begin
              reg308 <= "ZL9SEVIq9Z0ololHzi6D";
              reg309 <= $unsigned((($signed(reg304[(2'h3):(2'h2)]) ?
                  $signed("zNLOPEV") : ((7'h41) ?
                      (reg284 ^ reg311) : ((8'hac) ?
                          reg308 : reg276))) + ($unsigned(reg258[(4'ha):(3'h5)]) & "62ENGzdKFq63enWb")));
              reg310 <= forvar283[(4'he):(4'h9)];
            end
        end
    end
  module313 modinst350 (.y(wire349), .wire317(reg295), .wire315(forvar293), .wire316(reg308), .wire314(reg276), .clk(clk));
  assign wire351 = $signed($unsigned("chlH"));
  module352 modinst392 (wire391, clk, wire271, reg270, reg277, reg292, reg298);
  assign wire393 = (~&(~^($unsigned((reg252 ? reg303 : reg281)) ?
                       ((forvar287 > reg281) && (~|wire198)) : $signed((reg280 && reg290)))));
  always
    @(posedge clk) begin
      reg394 = {"DAWO",
          ({((~&(8'hac)) >= (^~reg265)),
              (^(reg300 ? forvar253 : (8'ha3)))} < {reg301[(3'h6):(1'h1)]})};
      for (forvar395 = (1'h0); (forvar395 < (1'h1)); forvar395 = (forvar395 + (1'h1)))
        begin
          reg396 <= "aMzMJZiiJrNxeQv";
        end
      reg397 = reg297;
      if ($unsigned($unsigned("lxAw3vrwLsRUsNSUPulgT")))
        begin
          for (forvar398 = (1'h0); (forvar398 < (1'h1)); forvar398 = (forvar398 + (1'h1)))
            begin
              reg399 = (-{forvar307, "oibr8DOQkOWSQ42n5"});
              reg400 <= "m2gwIt";
              reg401 <= {(8'h9e)};
            end
          if ((!(^reg256)))
            begin
              reg402 <= $signed(wire195);
            end
          else
            begin
              reg402 <= (forvar278[(3'h5):(1'h1)] + forvar287[(1'h1):(1'h0)]);
              reg403 <= {$unsigned((("AlCRtouTFwpHB" ?
                          {forvar278, reg270} : $signed(reg400)) ?
                      $signed(reg256[(3'h7):(3'h7)]) : reg252[(2'h2):(1'h1)])),
                  ((!wire251[(4'h8):(2'h2)]) ?
                      (^~($signed(reg312) == $unsigned(reg265))) : forvar293)};
              reg404 <= "S";
              reg405 <= ((reg296 ?
                  $signed(($signed(reg257) ?
                      $signed((8'hb3)) : wire197)) : (!$unsigned($signed(reg292)))) << (~|reg397[(1'h1):(1'h0)]));
              reg406 <= forvar287;
            end
          if (reg406[(1'h0):(1'h0)])
            begin
              reg407 <= ($unsigned($unsigned((!"g1hmk0p"))) ?
                  reg282 : "rN1AQQQh6cJzZMlTs0N");
              reg408 <= reg289;
            end
          else
            begin
              reg407 = $signed((|$unsigned("y")));
              reg408 <= (reg277[(1'h1):(1'h1)] ?
                  {($signed(reg258[(5'h14):(2'h2)]) > (~|$signed(reg394)))} : (("R0TT" ?
                          $signed((reg281 ?
                              (8'ha5) : reg301)) : $signed((reg304 >= reg299))) ?
                      (-forvar290[(4'hb):(4'ha)]) : reg309));
              reg409 <= (!"J8M2yYixsbZLW7cN");
              reg410 <= reg289[(4'h8):(3'h7)];
            end
          reg411 <= $unsigned({reg308, ((&"TUuZphQkV2ERvVnnRIP") ^~ reg260)});
        end
      else
        begin
          for (forvar398 = (1'h0); (forvar398 < (1'h1)); forvar398 = (forvar398 + (1'h1)))
            begin
              reg399 <= (~&"0XYFBUK");
            end
          for (forvar400 = (1'h0); (forvar400 < (3'h4)); forvar400 = (forvar400 + (1'h1)))
            begin
              reg401 <= ((!{(~^(&wire251))}) ?
                  {$signed((|(wire198 ? forvar278 : (8'hae)))),
                      ((7'h48) >= reg400)} : reg399[(4'hf):(4'he)]);
            end
          reg402 <= (($unsigned($unsigned($unsigned((8'hab)))) ?
              $unsigned(reg265[(1'h0):(1'h0)]) : "X6zJdy1g7") && "zrY6DTvnuXcHBFCw2miMPn");
          reg403 = "Alg4N19G9p7HSXaEJqz";
        end
    end
  always
    @(posedge clk) begin
      for (forvar412 = (1'h0); (forvar412 < (2'h3)); forvar412 = (forvar412 + (1'h1)))
        begin
          if (reg396[(3'h4):(2'h2)])
            begin
              reg413 <= ((wire198 + "5bFIsv") == reg254);
              reg414 = reg405[(2'h3):(1'h1)];
            end
          else
            begin
              reg413 <= reg268;
              reg414 <= forvar395;
              reg415 <= $unsigned(($unsigned((-"KoyleUrd")) <<< ($signed("Ss5efq1M5KV7apHgU4oi3c") * wire351[(3'h7):(3'h7)])));
              reg416 <= $unsigned((8'hb9));
            end
          if ("fh")
            begin
              reg417 <= $signed((~^"kQuFHbB4z3nqP"));
              reg418 <= $unsigned($signed(($signed(reg312) + $signed((reg259 || reg269)))));
              reg419 <= "1RAtqCWqSKqXy";
            end
          else
            begin
              reg417 <= forvar253[(4'h9):(4'h8)];
              reg418 <= "OHM2QoGbvapRJc57q7Am";
              reg419 <= wire349[(4'h9):(4'h9)];
              reg420 <= wire249;
            end
          reg421 <= (((^~reg265) && reg257) * $signed({reg411}));
          for (forvar422 = (1'h0); (forvar422 < (1'h1)); forvar422 = (forvar422 + (1'h1)))
            begin
              reg423 <= forvar253;
              reg424 <= {$signed((reg260[(3'h4):(1'h0)] ?
                      (^$unsigned((8'hae))) : "ze0MNB")),
                  ("om9LKHkD13y7TEh" ?
                      (({reg306, reg267} >> (~^forvar290)) ^~ $signed((wire251 ?
                          wire273 : reg256))) : reg258)};
              reg425 <= wire349[(2'h3):(2'h2)];
              reg426 <= forvar266;
            end
          reg427 <= ("N06Q2A2DIN0kTT2L1G5fT9" ?
              $unsigned($unsigned(forvar398)) : reg308[(4'ha):(2'h2)]);
        end
      for (forvar428 = (1'h0); (forvar428 < (3'h4)); forvar428 = (forvar428 + (1'h1)))
        begin
          if (($signed(reg419) ? (&"IEVM8EHIeCFRPX8") : $unsigned(reg415)))
            begin
              reg429 = $signed($signed("7dM7llyALc"));
            end
          else
            begin
              reg429 <= ($signed(((~^reg290[(4'hf):(4'hc)]) ?
                      ("PTH4fy94TkeweQb2moFqq" ?
                          (reg404 ? reg298 : reg285) : {reg276,
                              reg425}) : reg256[(2'h3):(1'h1)])) ?
                  $signed("PhUnaJwJI9Jv6o4") : ("yQzdrG" ?
                      ("04" ~^ reg300) : ((~|(reg303 ? wire251 : forvar274)) ?
                          ({(8'hb2)} ?
                              $unsigned((7'h48)) : $unsigned(reg268)) : ($unsigned(reg276) == reg411))));
            end
          reg430 <= $signed($signed("HLFUfMhLR62pJFgc7i"));
          for (forvar431 = (1'h0); (forvar431 < (2'h2)); forvar431 = (forvar431 + (1'h1)))
            begin
              reg432 <= (((($signed(reg280) ?
                      (!reg302) : reg287[(5'h15):(4'hc)]) && (~^(reg303 ?
                      reg304 : reg400))) - "xVnF1f") ?
                  "GyAG9CwvVXz" : {("0D" ?
                          $signed((wire271 ^~ reg430)) : "35iHPvqzv7FWzBBZsI6")});
              reg433 <= $unsigned((|reg258));
              reg434 <= reg278[(4'hc):(2'h3)];
            end
          reg435 <= ((({$signed((8'h9c)),
              (+reg403)} << "iwJZb") >>> reg300[(3'h6):(2'h3)]) ^~ ($unsigned(((|reg286) >>> (reg276 ?
              reg302 : (7'h41)))) <<< $signed("LDFKe7mQRkqwvIMsQGLPMS")));
        end
    end
  assign wire436 = "rKIPvdJuXV0XhxEcM0XYr";
  assign wire437 = ({(-(!(wire436 & (8'hb7))))} * $signed(($signed((reg259 ?
                       reg311 : reg423)) ~^ reg423)));
  module438 modinst519 (wire518, clk, forvar266, reg282, reg303, reg308, forvar253);
  always
    @(posedge clk) begin
      if (({reg434, $unsigned($unsigned($signed(reg426)))} ?
          reg308[(3'h6):(1'h0)] : $unsigned("")))
        begin
          reg520 <= reg277;
          if ((8'hb6))
            begin
              reg521 <= "ON64518uUt0";
            end
          else
            begin
              reg521 <= $signed(("a0QL7J4aUvMqf3" ?
                  reg255[(3'h5):(1'h1)] : $unsigned({(8'h9e)})));
              reg522 <= $signed(("5POpEBTEmRfkaMhvki" <<< ($signed(reg423[(1'h0):(1'h0)]) ?
                  "MyOfkr" : $unsigned((reg429 ? reg296 : reg304)))));
              reg523 <= $signed($signed($signed(reg261[(2'h3):(2'h3)])));
            end
          reg524 <= $unsigned("");
        end
      else
        begin
          reg520 <= $signed(($unsigned("r2fs7aF") >>> {($unsigned(forvar422) >> (reg275 ?
                  (8'ha4) : forvar253))}));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module47
#(parameter param153 = (&(~|(8'hbc))))
(y, clk, wire52, wire51, wire50, wire49, wire48);
  output wire [(32'h552):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'ha):(1'h0)] wire52;
  input wire signed [(4'hf):(1'h0)] wire51;
  input wire signed [(5'h12):(1'h0)] wire50;
  input wire signed [(5'h17):(1'h0)] wire49;
  input wire [(5'h12):(1'h0)] wire48;
  wire signed [(2'h2):(1'h0)] wire152;
  reg [(5'h14):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg150 = (1'h0);
  reg [(4'h8):(1'h0)] forvar149 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg146 = (1'h0);
  reg signed [(4'he):(1'h0)] reg145 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg144 = (1'h0);
  reg [(4'hf):(1'h0)] forvar143 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg142 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg141 = (1'h0);
  reg [(3'h5):(1'h0)] reg140 = (1'h0);
  reg [(2'h3):(1'h0)] reg139 = (1'h0);
  reg [(2'h3):(1'h0)] forvar138 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg137 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg136 = (1'h0);
  wire [(5'h10):(1'h0)] wire135;
  wire [(5'h12):(1'h0)] wire134;
  wire [(4'hd):(1'h0)] wire133;
  wire signed [(4'ha):(1'h0)] wire132;
  wire [(3'h4):(1'h0)] wire131;
  wire signed [(3'h6):(1'h0)] wire130;
  wire [(5'h15):(1'h0)] wire129;
  reg signed [(5'h16):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg122 = (1'h0);
  reg [(4'hc):(1'h0)] reg119 = (1'h0);
  reg [(4'h9):(1'h0)] forvar115 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg113 = (1'h0);
  reg [(4'hc):(1'h0)] reg127 = (1'h0);
  reg signed [(4'he):(1'h0)] reg126 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg125 = (1'h0);
  reg [(4'ha):(1'h0)] reg124 = (1'h0);
  reg [(4'he):(1'h0)] reg123 = (1'h0);
  reg [(5'h15):(1'h0)] forvar122 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg121 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg120 = (1'h0);
  reg [(3'h7):(1'h0)] forvar119 = (1'h0);
  reg signed [(4'he):(1'h0)] reg118 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg117 = (1'h0);
  reg [(5'h13):(1'h0)] reg116 = (1'h0);
  reg [(5'h11):(1'h0)] reg115 = (1'h0);
  reg [(5'h16):(1'h0)] reg114 = (1'h0);
  reg [(3'h7):(1'h0)] forvar113 = (1'h0);
  reg [(4'hc):(1'h0)] reg112 = (1'h0);
  reg [(3'h5):(1'h0)] reg111 = (1'h0);
  reg [(5'h16):(1'h0)] reg110 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg108 = (1'h0);
  reg [(3'h4):(1'h0)] forvar107 = (1'h0);
  reg [(5'h11):(1'h0)] reg106 = (1'h0);
  reg [(3'h7):(1'h0)] reg105 = (1'h0);
  reg [(4'hb):(1'h0)] forvar104 = (1'h0);
  reg [(4'hf):(1'h0)] reg103 = (1'h0);
  reg signed [(4'he):(1'h0)] reg101 = (1'h0);
  reg [(5'h11):(1'h0)] reg102 = (1'h0);
  reg [(3'h6):(1'h0)] forvar101 = (1'h0);
  reg [(4'h9):(1'h0)] reg100 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg99 = (1'h0);
  reg [(2'h2):(1'h0)] reg98 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar97 = (1'h0);
  reg [(5'h15):(1'h0)] reg96 = (1'h0);
  reg [(5'h16):(1'h0)] reg95 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg94 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar92 = (1'h0);
  reg signed [(4'he):(1'h0)] reg91 = (1'h0);
  reg [(2'h2):(1'h0)] reg90 = (1'h0);
  reg [(5'h13):(1'h0)] reg89 = (1'h0);
  reg [(5'h15):(1'h0)] reg88 = (1'h0);
  reg [(5'h16):(1'h0)] reg87 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg86 = (1'h0);
  reg [(5'h13):(1'h0)] reg85 = (1'h0);
  reg signed [(4'he):(1'h0)] reg84 = (1'h0);
  reg [(4'hd):(1'h0)] reg83 = (1'h0);
  reg [(5'h10):(1'h0)] reg82 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg81 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar80 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg79 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg78 = (1'h0);
  reg [(4'hb):(1'h0)] reg77 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg76 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg75 = (1'h0);
  reg [(4'hb):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg73 = (1'h0);
  reg [(5'h11):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg72 = (1'h0);
  reg [(5'h12):(1'h0)] forvar71 = (1'h0);
  reg [(5'h11):(1'h0)] reg70 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg69 = (1'h0);
  reg [(4'hc):(1'h0)] reg68 = (1'h0);
  reg [(4'hd):(1'h0)] reg67 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg66 = (1'h0);
  reg [(5'h13):(1'h0)] reg65 = (1'h0);
  reg [(5'h17):(1'h0)] reg61 = (1'h0);
  reg [(4'h9):(1'h0)] forvar54 = (1'h0);
  reg [(2'h3):(1'h0)] reg64 = (1'h0);
  reg [(3'h4):(1'h0)] reg63 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar61 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg60 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg59 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg58 = (1'h0);
  reg [(2'h3):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg56 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg55 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg54 = (1'h0);
  wire [(4'hc):(1'h0)] wire53;
  assign y = {wire152,
                 reg151,
                 reg150,
                 forvar149,
                 reg148,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 forvar143,
                 reg142,
                 reg141,
                 reg140,
                 reg139,
                 forvar138,
                 reg137,
                 reg136,
                 wire135,
                 wire134,
                 wire133,
                 wire132,
                 wire131,
                 wire130,
                 wire129,
                 reg128,
                 reg122,
                 reg119,
                 forvar115,
                 reg113,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 forvar122,
                 reg121,
                 reg120,
                 forvar119,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 forvar113,
                 reg112,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 forvar107,
                 reg106,
                 reg105,
                 forvar104,
                 reg103,
                 reg101,
                 reg102,
                 forvar101,
                 reg100,
                 reg99,
                 reg98,
                 forvar97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 forvar92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 forvar80,
                 reg79,
                 reg78,
                 reg77,
                 reg76,
                 reg75,
                 reg74,
                 reg73,
                 reg71,
                 reg72,
                 forvar71,
                 reg70,
                 reg69,
                 reg68,
                 reg67,
                 reg66,
                 reg65,
                 reg61,
                 forvar54,
                 reg64,
                 reg63,
                 reg62,
                 forvar61,
                 reg60,
                 reg59,
                 reg58,
                 reg57,
                 reg56,
                 reg55,
                 reg54,
                 wire53,
                 (1'h0)};
  assign wire53 = {wire49, $unsigned(wire52[(4'h9):(3'h7)])};
  always
    @(posedge clk) begin
      if ($unsigned(wire49[(5'h13):(4'h9)]))
        begin
          if ((($unsigned($unsigned((!(8'ha5)))) ?
              "FECXRckf7l9JwqPFY1Vm" : ("k" ?
                  $unsigned((+wire52)) : (+(-wire48)))) >= ("iaACaF1qygCaRDx" ?
              $signed((|"sLBBqhZTwADrEkIYAiwity")) : ((((7'h46) != wire53) ?
                  "3kSJaROn1N3xGFzSuZ08mq" : $unsigned(wire48)) >>> (wire48[(4'hf):(3'h7)] ?
                  wire50[(4'ha):(3'h6)] : "iLouAg5h2FQ4QcG7")))))
            begin
              reg54 = wire50;
            end
          else
            begin
              reg54 <= wire48;
            end
          reg55 = $unsigned(wire49);
          reg56 <= (reg55[(2'h2):(2'h2)] | $signed(($unsigned($signed(wire51)) ?
              wire51 : wire53)));
          if ((&$unsigned($signed(($unsigned(wire52) ?
              wire53 : $unsigned(reg55))))))
            begin
              reg57 <= wire52[(3'h5):(3'h4)];
              reg58 <= reg54;
              reg59 = $unsigned($unsigned((wire49[(2'h2):(2'h2)] < (~^$signed(reg57)))));
              reg60 <= (reg57[(1'h0):(1'h0)] & reg59);
            end
          else
            begin
              reg57 <= reg56[(4'hf):(3'h5)];
              reg58 <= ({$unsigned(({(8'hb7)} ?
                      $unsigned(reg54) : $unsigned(wire48))),
                  (($unsigned(wire51) ?
                          "885A0maHMLn0twI6b0qi" : wire49[(4'hb):(3'h4)]) ?
                      "iQ" : ($unsigned(reg56) ?
                          reg57 : ((7'h44) ?
                              reg57 : reg56)))} - ("SNxXwPCiXWWWhOA5uHk3" & (7'h41)));
              reg59 <= ($unsigned(reg56[(5'h11):(5'h11)]) ?
                  "XYNqRwRktR9pzpMtk" : (($signed((reg56 * wire51)) ?
                          $signed((~^wire48)) : $signed($signed(reg57))) ?
                      (~^"UCYPX") : (&wire48[(4'hf):(4'hc)])));
            end
          for (forvar61 = (1'h0); (forvar61 < (3'h4)); forvar61 = (forvar61 + (1'h1)))
            begin
              reg62 <= (~$signed((^(^{wire50, wire48}))));
              reg63 = (forvar61 ?
                  ("6HnwtA" ^ $unsigned(((!reg55) ?
                      reg60 : $signed(wire49)))) : "");
              reg64 = $unsigned($signed(forvar61));
            end
        end
      else
        begin
          for (forvar54 = (1'h0); (forvar54 < (2'h3)); forvar54 = (forvar54 + (1'h1)))
            begin
              reg55 <= (~^((((reg64 == reg56) ?
                      "GH4lE3lywxaWEOUe" : $unsigned(forvar54)) ?
                  $unsigned(reg55[(1'h0):(1'h0)]) : wire48) == reg63));
              reg56 = (reg64 ?
                  reg64[(1'h1):(1'h1)] : $unsigned((reg60[(2'h3):(2'h3)] ?
                      (+wire52) : reg57[(1'h0):(1'h0)])));
              reg57 <= wire50;
              reg58 <= (8'hb4);
              reg59 <= (+(~&(~^$signed((reg60 ? reg60 : reg59)))));
            end
          if ((|(8'hbc)))
            begin
              reg60 = wire48;
              reg61 <= (!wire48);
            end
          else
            begin
              reg60 <= "wfsBqO3sLdCW";
              reg61 <= ("" < reg56[(5'h12):(1'h0)]);
              reg62 = reg61[(2'h2):(2'h2)];
            end
          if (reg62)
            begin
              reg63 <= $signed(((reg56[(3'h7):(1'h0)] <= {(reg54 ?
                      wire51 : (7'h41))}) & (^~(~^((8'ha1) ?
                  reg59 : wire50)))));
              reg64 <= (|($signed($unsigned((wire53 < reg62))) ^ "857a"));
              reg65 <= ($unsigned(((+(reg60 ?
                      reg55 : (8'hb1))) < (wire53 + forvar54))) ?
                  wire51[(1'h1):(1'h1)] : wire50);
              reg66 <= (^~wire52);
            end
          else
            begin
              reg63 <= "W";
              reg64 <= ((+"Sz71v61q8uK9r6izHqD") ?
                  "W0Z2PruF8gI" : "m0lzYHonga");
              reg65 = $unsigned((^reg62));
              reg66 <= ("cEanxGG8sk4qO" ~^ "pmgDhfpUS1kJebAPeuJFBN");
            end
          reg67 <= (&$signed((+(reg65[(5'h11):(4'ha)] - reg62[(5'h12):(4'h9)]))));
          reg68 <= ((~$unsigned($signed((forvar61 ?
              reg61 : reg59)))) >> "dFEXqPPaY");
        end
      reg69 <= reg68[(4'h9):(4'h9)];
      if ("F4RuxNemekMEQz504")
        begin
          reg70 <= {$signed((~((forvar61 ?
                  reg61 : wire51) ^~ ((8'ha5) ^~ reg54)))),
              reg56};
          for (forvar71 = (1'h0); (forvar71 < (2'h3)); forvar71 = (forvar71 + (1'h1)))
            begin
              reg72 <= ({$signed(reg61[(2'h3):(1'h0)]),
                  "L65PuKi"} < (($unsigned((wire52 - (8'hb4))) << reg57) ?
                  reg70 : (({reg69, forvar54} || (reg70 ?
                      (7'h44) : (7'h45))) <<< ((^~reg67) ^ $unsigned(reg62)))));
            end
        end
      else
        begin
          if ((($signed("ItbTHfgb6h0VoMa8SHz") & "5nTCqx7W") & reg70))
            begin
              reg70 <= ((8'had) ?
                  $unsigned("tdwaL3gEUpAHQdkCWGGK8") : "Ylgthfy4xkHUaJl");
              reg71 <= reg68[(2'h2):(2'h2)];
              reg72 <= $unsigned($signed(((8'hbd) ?
                  "plk8" : $signed((wire50 ? reg59 : reg54)))));
              reg73 = ("PPo" ?
                  $signed((reg65[(4'hf):(2'h2)] ?
                      $unsigned((|reg71)) : $signed((reg56 | (7'h43))))) : reg56);
              reg74 <= "zop8rpN";
            end
          else
            begin
              reg70 <= {(("rs2q5hFQyXB" ? "sWYEWb2oC2S5013BBIouSO" : "e") ?
                      ((&reg73) <<< ((+reg60) ?
                          (forvar71 ~^ reg72) : reg69)) : "")};
              reg71 <= (forvar71[(4'h8):(1'h0)] - (^~("Gl20rYB7PiRhFONYc" << reg60)));
              reg72 <= {$signed(wire50)};
            end
          if ({({{reg57, (reg55 && reg69)}, $unsigned("pUzFx65Wu")} ?
                  wire51 : "Q")})
            begin
              reg75 <= (|(~|(~^$signed((^~reg64)))));
            end
          else
            begin
              reg75 <= $signed(("CFJE" || reg61[(1'h1):(1'h0)]));
              reg76 <= wire50;
              reg77 <= ((~&$signed(reg73[(2'h3):(2'h3)])) <= wire50[(2'h3):(2'h2)]);
              reg78 <= reg71;
              reg79 <= wire51;
            end
          for (forvar80 = (1'h0); (forvar80 < (2'h3)); forvar80 = (forvar80 + (1'h1)))
            begin
              reg81 = wire50[(3'h5):(1'h0)];
              reg82 <= reg67[(3'h4):(2'h3)];
              reg83 = reg78;
              reg84 <= (~^($unsigned((^{reg72, reg82})) ?
                  $unsigned($signed(forvar54[(2'h3):(1'h0)])) : reg72));
            end
          if (($unsigned((reg68 + ((wire51 ? reg54 : reg70) ?
              ((8'hbc) ~^ reg63) : (reg55 ? wire51 : (7'h48))))) << (((~|{reg69,
                  wire49}) != wire48[(5'h11):(4'hd)]) ?
              (~^(^~$unsigned(reg65))) : "5VZx3T1dk")))
            begin
              reg85 = ((8'hba) ?
                  "mJ51lvydaRUB2a" : ("7Pqp" ?
                      $unsigned(reg56[(1'h0):(1'h0)]) : (forvar61 == (|(~&wire52)))));
              reg86 <= "lZoar8hJZhHl5ibAK3";
            end
          else
            begin
              reg85 <= (($signed("XU9vfdgICQtKfiVNU8L61u") ?
                      $unsigned({(reg82 >= wire52),
                          (reg60 ? reg64 : wire51)}) : $signed((((8'h9e) ?
                          reg71 : reg56) & (reg77 ? reg62 : reg56)))) ?
                  $unsigned((reg84[(2'h2):(1'h1)] < ((reg75 ?
                          reg85 : forvar80) ?
                      wire49 : $unsigned(reg77)))) : (reg64[(1'h0):(1'h0)] ?
                      (~("S5uV" ?
                          "rkEqB2YYs" : ((8'ha3) << wire48))) : $signed(reg79)));
              reg86 <= ("geqrVbVEgk5NSnWtV4" ? reg63 : (|reg58[(3'h4):(1'h1)]));
              reg87 <= (&((reg82[(4'hb):(3'h5)] != reg83) ?
                  $signed(wire51) : $unsigned({$unsigned((7'h44)),
                      "VA2MoXg9XMbHMgmx6"})));
              reg88 <= forvar61[(4'h8):(1'h0)];
            end
          if (((reg86 ?
              $signed($signed("Q92ZW1w0mdwGO")) : ($signed("9U6zpOtid") ?
                  ($unsigned(reg79) * $signed(reg78)) : reg75)) >>> "yfEUgd"))
            begin
              reg89 <= "Dq";
              reg90 <= reg73[(2'h3):(1'h1)];
            end
          else
            begin
              reg89 <= $unsigned(reg74[(1'h1):(1'h1)]);
              reg90 <= (reg76[(4'hb):(4'hb)] && ($signed(((|reg57) >>> {reg86,
                      (8'hb4)})) ?
                  ({(reg55 <= reg84)} ?
                      $unsigned({reg89,
                          reg63}) : reg69[(2'h3):(1'h0)]) : (~{reg73})));
              reg91 <= {{$signed(reg60[(1'h0):(1'h0)])}, wire53};
            end
        end
    end
  always
    @(posedge clk) begin
      if (reg54[(3'h5):(3'h4)])
        begin
          for (forvar92 = (1'h0); (forvar92 < (2'h2)); forvar92 = (forvar92 + (1'h1)))
            begin
              reg93 <= ($unsigned($signed($unsigned($unsigned(reg85)))) ~^ reg64);
              reg94 <= ({reg79,
                      ((&reg87[(4'he):(2'h2)]) ?
                          "wpsKwg5Sz0danNkOPR" : $signed($signed(reg57)))} ?
                  $unsigned(reg61) : ($signed("JfTfc9skYrPOdNFW4oaOO") ?
                      ((reg73 ? (~forvar71) : ((8'ha4) ? reg69 : wire48)) ?
                          $unsigned($signed(reg59)) : $unsigned($unsigned(forvar92))) : (!((|(8'hb9)) << (|reg85)))));
              reg95 <= ($signed($unsigned((reg72 >= $signed(reg91)))) | forvar61[(2'h3):(2'h3)]);
            end
          reg96 <= $unsigned($signed({reg56, reg61}));
          for (forvar97 = (1'h0); (forvar97 < (1'h1)); forvar97 = (forvar97 + (1'h1)))
            begin
              reg98 <= {(-((^~wire51[(3'h5):(3'h4)]) ?
                      "cJY2qGXfc4P5snF" : ((wire53 ? (8'ha6) : reg91) ?
                          (reg81 ? reg87 : reg55) : "tiLEd"))),
                  ((((reg84 << (7'h48)) ?
                          "zTXFx1A9M4nyIEUp72fA" : $signed(reg96)) ?
                      $unsigned($signed(reg91)) : "rIqK") ~^ reg63[(1'h1):(1'h1)])};
            end
          reg99 <= ($unsigned("mGd9zbxb1yxOPCa1m") ?
              {{$signed($unsigned(reg54))}} : $signed(reg59[(4'ha):(3'h6)]));
          reg100 <= "yp2RNPc4yqA";
        end
      else
        begin
          for (forvar92 = (1'h0); (forvar92 < (2'h3)); forvar92 = (forvar92 + (1'h1)))
            begin
              reg93 <= "XBCSQiPIvdIucLZZAIBf";
              reg94 <= $unsigned((reg72[(1'h0):(1'h0)] | ((reg84 ?
                      (forvar71 ? reg86 : reg90) : (reg89 ? reg95 : reg75)) ?
                  "RTAfdSrqcGQRai5ihf5oQq" : reg88)));
            end
          reg95 <= (((~|({reg82, forvar92} ?
                  (&reg59) : (reg72 != (8'hae)))) != "o81qpHoeh4ofgM") ?
              reg64 : (+(~|reg59)));
        end
      if ("uhWQusT")
        begin
          for (forvar101 = (1'h0); (forvar101 < (1'h1)); forvar101 = (forvar101 + (1'h1)))
            begin
              reg102 <= $unsigned($signed($signed(({reg85} ?
                  (~^(8'haf)) : "ZXpiGNgs8yIgPRatVL4"))));
            end
        end
      else
        begin
          if ($unsigned($unsigned(reg76)))
            begin
              reg101 <= (8'ha0);
              reg102 <= $unsigned({((-$signed(wire51)) ?
                      $unsigned($signed(reg67)) : $signed("M2YwZKFrAh")),
                  {{((7'h41) ? reg54 : reg81), (^~wire48)}}});
              reg103 <= (reg66[(3'h6):(2'h3)] <= $signed((+("e3kvJd5ZdEcXtYnfnDa3" ^~ (reg89 <<< forvar80)))));
            end
          else
            begin
              reg101 <= ($signed(("AybdECh4fKvv8Teb" ?
                      ({(8'hb5),
                          reg64} - $signed((8'h9f))) : reg103[(4'h9):(4'h8)])) ?
                  (~&reg65[(4'ha):(1'h0)]) : reg65[(3'h5):(3'h5)]);
              reg102 <= "EgVYfObhHwppOQ2";
            end
          for (forvar104 = (1'h0); (forvar104 < (1'h0)); forvar104 = (forvar104 + (1'h1)))
            begin
              reg105 = (-$unsigned({$signed(reg100)}));
              reg106 <= reg61[(4'hc):(1'h0)];
            end
          for (forvar107 = (1'h0); (forvar107 < (2'h2)); forvar107 = (forvar107 + (1'h1)))
            begin
              reg108 <= (~|reg55);
              reg109 = $signed({reg77});
              reg110 <= (reg60 || "k");
              reg111 <= reg74[(4'ha):(3'h6)];
            end
        end
      reg112 = {(~^(|("roV8TEZvXSplMh7UrtTc" ?
              (reg87 ? (7'h40) : (8'hb8)) : (forvar80 < reg110))))};
      if ((forvar80[(1'h1):(1'h0)] || ($unsigned({forvar92[(3'h4):(1'h1)]}) ?
          {((!reg77) ? {reg81, reg88} : {reg86, (8'hbb)})} : (~&(~&forvar80)))))
        begin
          for (forvar113 = (1'h0); (forvar113 < (2'h3)); forvar113 = (forvar113 + (1'h1)))
            begin
              reg114 <= $signed($signed(($signed(forvar80) ^ ($unsigned(reg57) ~^ "xsyvhUyqhaqa"))));
              reg115 <= $signed(("" ?
                  reg59 : {{forvar92, ((8'hb9) + (8'hbe))},
                      $signed($unsigned(reg54))}));
              reg116 <= (^~$unsigned({reg99[(3'h6):(3'h5)],
                  $unsigned((reg114 && forvar97))}));
              reg117 <= "cNAFepJipaII";
              reg118 = "abX3";
            end
          for (forvar119 = (1'h0); (forvar119 < (2'h2)); forvar119 = (forvar119 + (1'h1)))
            begin
              reg120 <= ((~reg61[(4'hd):(4'h8)]) != (reg69[(2'h2):(1'h0)] ?
                  (+$unsigned(forvar54)) : forvar92[(2'h2):(1'h1)]));
              reg121 <= $signed(reg106);
            end
          for (forvar122 = (1'h0); (forvar122 < (2'h2)); forvar122 = (forvar122 + (1'h1)))
            begin
              reg123 <= $signed($signed(reg114[(5'h11):(3'h5)]));
              reg124 <= (8'ha7);
              reg125 <= ((reg109[(3'h7):(3'h7)] ?
                      {forvar92[(1'h0):(1'h0)]} : $signed($signed($unsigned((8'hac))))) ?
                  reg87[(4'he):(2'h3)] : {$signed($unsigned((reg124 ?
                          forvar54 : forvar97)))});
              reg126 <= reg77[(4'ha):(1'h0)];
              reg127 <= $unsigned(reg121[(3'h4):(2'h2)]);
            end
        end
      else
        begin
          if ((reg91 != forvar92))
            begin
              reg113 <= ($unsigned({("eJHVu5ty" ?
                      $unsigned(reg69) : forvar97[(1'h1):(1'h0)]),
                  reg100}) <= $unsigned(reg126));
              reg114 <= ($unsigned({"S52olF", $signed($unsigned((8'h9c)))}) ?
                  (~reg96[(2'h3):(2'h2)]) : {reg54, (&(8'ha3))});
            end
          else
            begin
              reg113 <= $unsigned("8HCYXnuMS5");
              reg114 <= "dIzDXOkysqVUlfROD3i08J";
            end
          for (forvar115 = (1'h0); (forvar115 < (1'h0)); forvar115 = (forvar115 + (1'h1)))
            begin
              reg116 = $signed(wire51);
              reg117 <= reg110;
              reg118 <= "43diwhPm";
              reg119 <= $signed((^~reg117[(3'h6):(3'h5)]));
            end
          if (($unsigned(($signed((~^reg84)) ?
              reg111[(1'h1):(1'h0)] : {reg57[(1'h1):(1'h0)],
                  (~reg114)})) >>> $unsigned(reg90[(2'h2):(2'h2)])))
            begin
              reg120 <= (8'h9f);
              reg121 <= (($signed({(|reg123)}) ?
                  ($signed((~|reg70)) && reg56) : $unsigned(($signed(reg63) <<< (7'h40)))) <<< ($signed("AQyFW1Isl") >>> {reg85[(5'h13):(4'h9)],
                  reg111}));
              reg122 <= (forvar104 ?
                  (-(~$unsigned("rB0VehlBR3P7B9"))) : $signed((reg75[(5'h10):(4'ha)] == ($unsigned(reg127) == (8'h9d)))));
              reg123 <= reg83[(1'h1):(1'h0)];
            end
          else
            begin
              reg120 <= reg72[(2'h2):(1'h1)];
              reg121 <= {$signed(forvar115)};
              reg122 = (wire48[(4'he):(3'h6)] ?
                  ("0G" < "rONhbGpKR3mEdUQJMO7") : {$unsigned($unsigned($unsigned(forvar104))),
                      (!("Nk4hW8Rrf633uAVxpF" >> reg59[(5'h16):(4'hf)]))});
            end
          reg124 = ($signed((|"8yK7uN")) + "urTlGTVaSbNJKueFVJ");
        end
    end
  always
    @(posedge clk) begin
      reg128 <= ($signed("6kKkIT8fxU1iiU") ? "nwMhfKJ" : reg78);
    end
  assign wire129 = (8'hbc);
  assign wire130 = $signed($signed(reg54[(3'h4):(3'h4)]));
  assign wire131 = {"3eFMXu8L8I4YTlWX"};
  assign wire132 = {$signed((reg125[(4'hb):(3'h4)] >> ((8'hba) ^ reg115))), ""};
  assign wire133 = {"an4Gzum"};
  assign wire134 = $signed((+wire53));
  assign wire135 = {reg95[(3'h6):(3'h6)], wire50};
  always
    @(posedge clk) begin
      reg136 <= (^"6yVZaYsywOSn5fQUlQTWn");
      reg137 <= (~&"bg5HYfAbIlSt");
      for (forvar138 = (1'h0); (forvar138 < (2'h3)); forvar138 = (forvar138 + (1'h1)))
        begin
          if ((+reg105[(2'h3):(2'h3)]))
            begin
              reg139 <= "5zIB";
              reg140 <= forvar119[(2'h3):(2'h3)];
              reg141 <= ((((8'h9c) >>> ((reg71 ? (7'h47) : reg122) - ((8'h9c) ?
                  reg94 : (8'h9e)))) ^ (("8aEZ9RR" >> $unsigned((8'ha8))) ?
                  "" : $unsigned("DAAibtYC"))) && (reg124[(1'h1):(1'h1)] ?
                  $unsigned(forvar80) : $signed(((^reg83) ?
                      ((8'ha9) > reg79) : (reg72 <<< reg55)))));
              reg142 <= $signed(wire130[(1'h1):(1'h0)]);
            end
          else
            begin
              reg139 <= $unsigned(((reg103 + reg77) ?
                  $unsigned(reg109) : $signed($unsigned({reg59}))));
              reg140 <= $unsigned(((~&reg102[(4'hb):(3'h7)]) && "ZS"));
            end
          for (forvar143 = (1'h0); (forvar143 < (1'h0)); forvar143 = (forvar143 + (1'h1)))
            begin
              reg144 <= (^($signed($signed((reg124 ? reg99 : (8'hb4)))) ?
                  "EDOvokGLw0LdvHREaTlgZ" : (reg95[(1'h1):(1'h0)] & ({reg54} <<< "WPYIJr1pJw1f2VCRTif"))));
              reg145 = $signed($unsigned(($unsigned((~&wire51)) ~^ {reg114})));
            end
          if ((({(~"8WdMecEdFHAUW3vFZfiO6i"),
                      ({(8'hb6), reg90} ?
                          (reg122 <<< reg96) : (reg71 ? (8'ha3) : reg66))} ?
                  $signed({((8'hbc) << reg109)}) : "WUqKkGOsP") ?
              (reg137[(3'h7):(3'h4)] || $unsigned(reg94[(3'h4):(1'h0)])) : $signed(reg121[(3'h4):(2'h2)])))
            begin
              reg146 <= reg55;
            end
          else
            begin
              reg146 <= ($signed(((&$unsigned(wire135)) >>> (reg103 ?
                      reg78[(3'h5):(1'h0)] : (~reg141)))) ?
                  (~|(^$signed({reg110, reg125}))) : (^~(reg84 ?
                      "m" : "KTF9qsFm7aZIkZ0")));
              reg147 <= {(&"Q8vqH")};
            end
          reg148 <= ((|reg73[(1'h0):(1'h0)]) ? forvar97 : reg78[(3'h6):(1'h1)]);
        end
      for (forvar149 = (1'h0); (forvar149 < (2'h2)); forvar149 = (forvar149 + (1'h1)))
        begin
          reg150 <= $unsigned($unsigned(($unsigned($signed(reg124)) != "1qoGyf")));
          reg151 <= $unsigned($signed($unsigned(reg126[(3'h7):(1'h0)])));
        end
    end
  assign wire152 = $unsigned("XOA86ZEQq6iSK64");
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module438  (y, clk, wire443, wire442, wire441, wire440, wire439);
  output wire [(32'h392):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire443;
  input wire signed [(5'h10):(1'h0)] wire442;
  input wire signed [(4'h9):(1'h0)] wire441;
  input wire signed [(4'hc):(1'h0)] wire440;
  input wire [(5'h17):(1'h0)] wire439;
  reg [(5'h10):(1'h0)] reg517 = (1'h0);
  reg [(5'h11):(1'h0)] reg516 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg515 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg514 = (1'h0);
  reg [(4'hc):(1'h0)] forvar513 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar512 = (1'h0);
  reg [(4'hc):(1'h0)] reg511 = (1'h0);
  reg [(5'h17):(1'h0)] reg510 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg509 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg508 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg507 = (1'h0);
  reg [(3'h4):(1'h0)] reg506 = (1'h0);
  reg [(2'h2):(1'h0)] forvar505 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar504 = (1'h0);
  wire [(2'h2):(1'h0)] wire503;
  wire signed [(4'he):(1'h0)] wire502;
  wire [(5'h16):(1'h0)] wire501;
  wire [(5'h16):(1'h0)] wire500;
  reg signed [(4'hb):(1'h0)] reg499 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg498 = (1'h0);
  reg [(4'hb):(1'h0)] reg497 = (1'h0);
  reg [(4'hc):(1'h0)] forvar496 = (1'h0);
  wire [(4'hb):(1'h0)] wire495;
  wire signed [(4'hc):(1'h0)] wire494;
  wire [(5'h14):(1'h0)] wire493;
  wire signed [(4'hf):(1'h0)] wire492;
  wire [(5'h11):(1'h0)] wire491;
  wire signed [(3'h7):(1'h0)] wire490;
  wire [(3'h5):(1'h0)] wire489;
  wire signed [(4'he):(1'h0)] wire488;
  wire signed [(5'h12):(1'h0)] wire487;
  wire signed [(3'h6):(1'h0)] wire486;
  reg signed [(3'h4):(1'h0)] reg485 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg484 = (1'h0);
  reg [(5'h13):(1'h0)] reg483 = (1'h0);
  reg signed [(4'he):(1'h0)] reg482 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg481 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar480 = (1'h0);
  reg [(5'h10):(1'h0)] reg479 = (1'h0);
  reg [(3'h5):(1'h0)] reg478 = (1'h0);
  reg [(5'h16):(1'h0)] reg477 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar476 = (1'h0);
  reg [(3'h6):(1'h0)] forvar475 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg474 = (1'h0);
  reg [(5'h15):(1'h0)] reg473 = (1'h0);
  reg [(4'hc):(1'h0)] reg472 = (1'h0);
  reg [(2'h2):(1'h0)] reg471 = (1'h0);
  reg [(3'h5):(1'h0)] reg470 = (1'h0);
  reg [(5'h16):(1'h0)] reg469 = (1'h0);
  reg [(3'h4):(1'h0)] reg468 = (1'h0);
  reg [(5'h13):(1'h0)] reg467 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar466 = (1'h0);
  reg [(4'ha):(1'h0)] reg465 = (1'h0);
  reg [(5'h12):(1'h0)] reg464 = (1'h0);
  reg [(4'he):(1'h0)] reg463 = (1'h0);
  reg [(3'h5):(1'h0)] forvar462 = (1'h0);
  reg [(4'hf):(1'h0)] forvar461 = (1'h0);
  reg [(3'h6):(1'h0)] reg460 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg459 = (1'h0);
  reg [(4'h9):(1'h0)] reg458 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg457 = (1'h0);
  reg [(5'h14):(1'h0)] reg456 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg455 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg454 = (1'h0);
  reg [(4'hc):(1'h0)] reg453 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg452 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg451 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg450 = (1'h0);
  reg [(3'h5):(1'h0)] reg449 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg448 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar447 = (1'h0);
  reg [(5'h13):(1'h0)] forvar446 = (1'h0);
  wire [(4'hc):(1'h0)] wire445;
  wire signed [(5'h10):(1'h0)] wire444;
  assign y = {reg517,
                 reg516,
                 reg515,
                 reg514,
                 forvar513,
                 forvar512,
                 reg511,
                 reg510,
                 reg509,
                 reg508,
                 reg507,
                 reg506,
                 forvar505,
                 forvar504,
                 wire503,
                 wire502,
                 wire501,
                 wire500,
                 reg499,
                 reg498,
                 reg497,
                 forvar496,
                 wire495,
                 wire494,
                 wire493,
                 wire492,
                 wire491,
                 wire490,
                 wire489,
                 wire488,
                 wire487,
                 wire486,
                 reg485,
                 reg484,
                 reg483,
                 reg482,
                 reg481,
                 forvar480,
                 reg479,
                 reg478,
                 reg477,
                 forvar476,
                 forvar475,
                 reg474,
                 reg473,
                 reg472,
                 reg471,
                 reg470,
                 reg469,
                 reg468,
                 reg467,
                 forvar466,
                 reg465,
                 reg464,
                 reg463,
                 forvar462,
                 forvar461,
                 reg460,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 reg454,
                 reg453,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 forvar447,
                 forvar446,
                 wire445,
                 wire444,
                 (1'h0)};
  assign wire444 = $signed({$signed(wire443), wire442[(1'h1):(1'h0)]});
  assign wire445 = wire439;
  always
    @(posedge clk) begin
      for (forvar446 = (1'h0); (forvar446 < (2'h3)); forvar446 = (forvar446 + (1'h1)))
        begin
          for (forvar447 = (1'h0); (forvar447 < (3'h4)); forvar447 = (forvar447 + (1'h1)))
            begin
              reg448 <= $signed((~$signed(wire440)));
              reg449 <= $unsigned(($unsigned({(wire439 + (8'hae))}) || $signed(wire441[(1'h1):(1'h1)])));
              reg450 <= (wire443 ?
                  (-forvar447[(2'h3):(2'h2)]) : $unsigned((8'hb7)));
            end
          if (({{$signed("5bgw")}} ?
              forvar446[(5'h11):(5'h10)] : forvar447[(4'h9):(1'h0)]))
            begin
              reg451 <= (+"Hodi747wFcF");
              reg452 <= wire444;
              reg453 = $unsigned($unsigned((^~"NeSxbYnTpworUYxik1z")));
            end
          else
            begin
              reg451 <= "ao";
              reg452 <= ((-wire443) ?
                  (($signed((^wire443)) != ((8'hae) <= "ou2FH")) ?
                      ((~^{wire445, wire445}) ?
                          "lfAQYChG2Id5lJi4NGX" : ($signed(reg449) ~^ (wire439 == wire445))) : wire444[(1'h0):(1'h0)]) : reg450[(3'h6):(1'h1)]);
              reg453 <= {reg452};
              reg454 <= (8'hb1);
              reg455 <= ((wire445[(4'ha):(2'h3)] >>> (-($unsigned(reg448) ?
                  (reg450 ? wire443 : wire444) : reg449))) << ("0w" ?
                  "qbwhScQzVkAvTiN5" : $unsigned({$signed(wire443), reg449})));
            end
          if ($signed(wire441))
            begin
              reg456 <= ((wire441[(3'h5):(3'h5)] ?
                      (+wire443) : ((7'h43) ~^ ($unsigned(wire445) ?
                          {wire443, reg450} : wire443))) ?
                  $signed("9JiQpbNSbKJ") : reg453);
              reg457 <= (+forvar447[(4'he):(3'h6)]);
              reg458 <= (($signed(reg456[(4'hc):(4'h9)]) && (^$signed($signed(reg451)))) | (("6QS0L" * (~|reg456)) != ((~reg448) ?
                  forvar446 : reg457[(1'h0):(1'h0)])));
              reg459 <= wire444[(3'h7):(2'h2)];
              reg460 <= ((wire443 + $unsigned({(8'ha8),
                  (reg456 ?
                      wire444 : (8'hb5))})) | $unsigned(wire445[(3'h5):(3'h4)]));
            end
          else
            begin
              reg456 = (((((8'ha3) ? reg449[(3'h4):(2'h3)] : (8'hba)) ?
                      ((wire440 || wire443) >>> reg457) : ("HgswDClZC9dL" ~^ "")) == (~($unsigned((8'hb0)) ^~ $unsigned(reg457)))) ?
                  (7'h41) : $unsigned($unsigned(((reg455 > reg449) ?
                      $signed(wire444) : (wire440 > wire439)))));
              reg457 = reg449[(1'h1):(1'h1)];
              reg458 <= wire439[(5'h14):(4'ha)];
              reg459 <= $unsigned(reg458);
            end
        end
      for (forvar461 = (1'h0); (forvar461 < (2'h3)); forvar461 = (forvar461 + (1'h1)))
        begin
          for (forvar462 = (1'h0); (forvar462 < (1'h1)); forvar462 = (forvar462 + (1'h1)))
            begin
              reg463 = (($unsigned(((forvar462 <<< reg450) ?
                  {(8'ha0), reg448} : {(8'hb0),
                      reg451})) <<< (^~{"4NBUz1zykp7F"})) + ((reg452 > ((forvar447 ?
                          reg457 : reg454) ?
                      (forvar447 >= reg452) : (7'h43))) ?
                  reg460[(3'h5):(1'h0)] : ((~{forvar446}) & {$signed(forvar447)})));
              reg464 <= ((|$signed($signed({forvar447}))) <= $unsigned(((~&reg455) ?
                  {"YRChWywbFl4OAqu4hvs",
                      (wire443 ? (8'h9d) : forvar462)} : "kgAse")));
            end
          reg465 = ($unsigned((~^(-wire442[(3'h5):(2'h3)]))) ?
              (reg448 != {((reg448 <= reg450) >= forvar462[(3'h5):(2'h2)])}) : (-$unsigned($unsigned(reg450))));
          for (forvar466 = (1'h0); (forvar466 < (1'h1)); forvar466 = (forvar466 + (1'h1)))
            begin
              reg467 <= reg463;
              reg468 = forvar461;
              reg469 = forvar446;
              reg470 <= ($signed(((^(reg465 ? reg450 : (8'hb4))) ?
                      ($signed(reg451) ?
                          (wire440 ?
                              wire443 : forvar462) : $unsigned((8'hba))) : "s")) ?
                  reg451[(2'h3):(1'h0)] : "1gnSKKOqmELaoSN");
            end
          reg471 <= wire441;
          if (($signed(wire442) ?
              {$signed(reg463[(4'hb):(3'h6)])} : $unsigned("0RLaxvSo8cAv")))
            begin
              reg472 <= $signed({{wire440[(2'h3):(1'h0)],
                      reg448[(3'h4):(2'h3)]},
                  $unsigned((!$unsigned(reg456)))});
            end
          else
            begin
              reg472 <= (~^$unsigned(reg465));
            end
        end
      reg473 <= (forvar446 ?
          "hATMKBWd3ry0RK" : (-{{(!reg455), $signed(reg469)},
              ((reg459 ? reg458 : wire441) ?
                  wire441[(4'h9):(4'h9)] : reg465[(4'h9):(3'h5)])}));
      reg474 <= $unsigned((|(reg448 ?
          (reg464 ?
              (forvar466 ^~ (8'haf)) : wire443) : ("H4JLvePGg8Pzd" >>> "f7tENwtx6vdtv3Dh"))));
      for (forvar475 = (1'h0); (forvar475 < (2'h2)); forvar475 = (forvar475 + (1'h1)))
        begin
          for (forvar476 = (1'h0); (forvar476 < (2'h3)); forvar476 = (forvar476 + (1'h1)))
            begin
              reg477 <= reg448[(3'h4):(2'h2)];
              reg478 = $unsigned(($signed(($unsigned((8'h9f)) ?
                  $unsigned(wire439) : reg454)) <<< ($unsigned((forvar447 ?
                      reg450 : reg460)) ?
                  $signed((forvar461 && reg468)) : $unsigned((^(8'h9e))))));
              reg479 <= reg474[(2'h3):(2'h2)];
            end
          for (forvar480 = (1'h0); (forvar480 < (2'h3)); forvar480 = (forvar480 + (1'h1)))
            begin
              reg481 <= $unsigned($signed((^~(wire440 ^ {reg456}))));
              reg482 = reg472;
              reg483 = ((~|{reg474,
                  (&(!wire443))}) - $unsigned(reg468[(1'h1):(1'h0)]));
              reg484 <= reg452[(2'h2):(1'h1)];
              reg485 <= ((!{(reg452[(3'h7):(3'h7)] ?
                      $signed(reg464) : "pd576R16elTfc")}) <<< (~^((~(reg456 ^ reg457)) << reg474)));
            end
        end
    end
  assign wire486 = $signed($signed((~&{(reg469 ? reg448 : forvar447),
                       {reg451}})));
  assign wire487 = ("9" <<< reg452);
  assign wire488 = "pKTRBs4J8G57B";
  assign wire489 = reg448;
  assign wire490 = reg469[(2'h3):(1'h1)];
  assign wire491 = (reg473 >= reg459[(4'hd):(4'hb)]);
  assign wire492 = reg460;
  assign wire493 = {$unsigned((7'h44))};
  assign wire494 = wire439;
  assign wire495 = wire491[(3'h7):(3'h5)];
  always
    @(posedge clk) begin
      for (forvar496 = (1'h0); (forvar496 < (2'h2)); forvar496 = (forvar496 + (1'h1)))
        begin
          reg497 <= "tO2gW0htqiCNkOni";
          reg498 <= $signed((8'ha7));
        end
      reg499 <= wire441[(3'h6):(1'h1)];
    end
  assign wire500 = (~&"qhL4u0Y7V26Ccq2pk");
  assign wire501 = $unsigned(reg465[(4'h9):(1'h1)]);
  assign wire502 = $unsigned($unsigned((&$unsigned((forvar480 ?
                       reg468 : reg457)))));
  assign wire503 = ({(-{{reg470,
                               reg456}})} <<< ($unsigned($unsigned("kY4pI")) + $signed($signed($signed(reg458)))));
  always
    @(posedge clk) begin
      for (forvar504 = (1'h0); (forvar504 < (3'h4)); forvar504 = (forvar504 + (1'h1)))
        begin
          for (forvar505 = (1'h0); (forvar505 < (2'h2)); forvar505 = (forvar505 + (1'h1)))
            begin
              reg506 <= $signed(wire503);
            end
          if ($unsigned(reg452[(4'h9):(3'h4)]))
            begin
              reg507 <= $signed($unsigned($unsigned((~|$unsigned((8'had))))));
              reg508 = ($signed({"R6oDzUpNqkwJ9",
                      ((reg499 ? forvar466 : reg478) ^~ (8'ha4))}) ?
                  "OFw" : "VFzID2k8");
              reg509 <= $signed(((~|((reg456 & wire439) ~^ $signed(wire439))) ?
                  wire444[(2'h2):(1'h1)] : $signed($signed((8'hb8)))));
              reg510 <= (-("YQpKF3V" ?
                  wire489[(1'h0):(1'h0)] : ($unsigned($signed(wire502)) + wire492[(1'h1):(1'h0)])));
              reg511 <= $signed("2f9Kqy");
            end
          else
            begin
              reg507 = ((~(!$signed($signed((8'haf))))) ?
                  $unsigned(((reg456[(3'h4):(2'h2)] ?
                      $unsigned(wire488) : (wire491 | (7'h41))) > reg455)) : reg455);
            end
        end
      for (forvar512 = (1'h0); (forvar512 < (2'h2)); forvar512 = (forvar512 + (1'h1)))
        begin
          for (forvar513 = (1'h0); (forvar513 < (2'h3)); forvar513 = (forvar513 + (1'h1)))
            begin
              reg514 <= "ZQUimnDn5H1U9";
              reg515 <= $signed((-"h6txJ"));
              reg516 = ($signed((("0oPWcyaQMrvhf" ?
                      "qB2IOgqEill0A1n1" : {reg515, wire503}) ?
                  ("xy5pWmaJq27HCFinJAV" > (reg458 <= wire487)) : ($unsigned(reg507) != $unsigned(reg470)))) << $signed((((wire500 ^~ (8'ha8)) ?
                      (wire503 ? (8'hac) : (8'ha6)) : (reg508 & forvar475)) ?
                  "v0w0yghBUu5RIeT7no" : "mH5FuEqWUz1lNYbX7x")));
              reg517 <= (reg514[(2'h2):(2'h2)] ?
                  (&(~|($unsigned(reg510) - $signed(reg507)))) : {$signed(forvar475)});
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module352
#( parameter param389 = (((!(((8'hb7) ? (8'hb0) : (8'ha2)) ? (+(8'hb2)) : ((7'h44) ? (8'hb7) : (8'hb6)))) ? {(((8'ha9) ? (8'ha4) : (8'ha2)) > (&(8'h9c)))} : (|(|((7'h40) ? (7'h41) : (8'hb5))))) >>> {((((8'ha4) ? (7'h46) : (8'ha0)) ? (~&(8'ha7)) : ((8'hb0) ? (8'hba) : (8'hb9))) ? (((8'hbe) || (8'hbf)) ~^ ((7'h46) ? (7'h44) : (8'hb1))) : (|((8'hae) ? (7'h48) : (8'had)))), (({(8'hab), (8'hb4)} ~^ {(8'hac)}) < (~&((8'ha0) ? (8'h9f) : (7'h41))))})
, parameter param390 = (((-(~^{(8'hb5), param389})) ? ({param389} ? ((~param389) ? param389 : ((8'ha5) - param389)) : (8'hb8)) : param389) ? param389 : ({((param389 ? param389 : param389) != (!param389))} <<< param389)) )
(y, clk, wire357, wire356, wire355, wire354, wire353);
  output wire [(32'h177):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire357;
  input wire signed [(4'hb):(1'h0)] wire356;
  input wire signed [(2'h3):(1'h0)] wire355;
  input wire [(2'h2):(1'h0)] wire354;
  input wire signed [(3'h7):(1'h0)] wire353;
  reg [(4'h9):(1'h0)] reg388 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg387 = (1'h0);
  wire [(2'h3):(1'h0)] wire386;
  wire [(4'h9):(1'h0)] wire385;
  wire [(5'h14):(1'h0)] wire384;
  wire [(5'h17):(1'h0)] wire383;
  wire signed [(4'h8):(1'h0)] wire382;
  wire [(3'h5):(1'h0)] wire381;
  wire signed [(4'ha):(1'h0)] wire380;
  wire [(5'h15):(1'h0)] wire379;
  wire signed [(4'hf):(1'h0)] wire378;
  wire signed [(5'h15):(1'h0)] wire377;
  wire [(3'h5):(1'h0)] wire376;
  reg [(3'h4):(1'h0)] reg375 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg374 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg373 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar372 = (1'h0);
  wire [(3'h7):(1'h0)] wire371;
  wire [(4'hc):(1'h0)] wire370;
  wire signed [(4'hf):(1'h0)] wire369;
  wire [(5'h13):(1'h0)] wire368;
  wire [(4'h9):(1'h0)] wire367;
  wire [(5'h11):(1'h0)] wire366;
  reg [(4'hf):(1'h0)] reg365 = (1'h0);
  reg [(3'h4):(1'h0)] forvar362 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg364 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg363 = (1'h0);
  reg [(5'h15):(1'h0)] reg362 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg361 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg360 = (1'h0);
  wire signed [(5'h15):(1'h0)] wire359;
  reg signed [(4'hd):(1'h0)] reg358 = (1'h0);
  assign y = {reg388,
                 reg387,
                 wire386,
                 wire385,
                 wire384,
                 wire383,
                 wire382,
                 wire381,
                 wire380,
                 wire379,
                 wire378,
                 wire377,
                 wire376,
                 reg375,
                 reg374,
                 reg373,
                 forvar372,
                 wire371,
                 wire370,
                 wire369,
                 wire368,
                 wire367,
                 wire366,
                 reg365,
                 forvar362,
                 reg364,
                 reg363,
                 reg362,
                 reg361,
                 reg360,
                 wire359,
                 reg358,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg358 <= {(&((^~(wire354 | wire354)) != wire357))};
    end
  assign wire359 = wire354;
  always
    @(posedge clk) begin
      if (wire355)
        begin
          if (("FQ" != ((|wire353) ?
              (wire359 + $unsigned(wire355)) : (&reg358[(4'h9):(1'h0)]))))
            begin
              reg360 <= {$unsigned((wire354 ?
                      wire354[(2'h2):(1'h1)] : $unsigned($signed(wire353))))};
            end
          else
            begin
              reg360 <= {(reg358 ?
                      $signed($signed(wire356)) : $signed($signed(wire357))),
                  ("4Vot39P89TG0" == $unsigned((~$signed(wire359))))};
              reg361 <= (wire356[(3'h5):(3'h5)] ?
                  {((8'hb4) & (7'h43)),
                      $unsigned($unsigned({(8'hb2)}))} : (reg360 ?
                      $signed({wire355[(2'h3):(1'h1)],
                          reg358[(1'h0):(1'h0)]}) : $unsigned($signed($signed(wire357)))));
              reg362 <= "Of8OcuU38cxNOpOh5";
              reg363 <= wire354[(1'h1):(1'h0)];
              reg364 = "9CtW4arB5c";
            end
        end
      else
        begin
          reg360 <= $signed((reg362[(4'hf):(4'hb)] ?
              $signed($signed({reg358})) : ((&"Q8CMHV0f1JquoY") > $unsigned((wire353 ?
                  reg358 : reg363)))));
          reg361 <= (($signed("FbVCMn") ~^ $signed((8'hbe))) | (7'h45));
          for (forvar362 = (1'h0); (forvar362 < (1'h1)); forvar362 = (forvar362 + (1'h1)))
            begin
              reg363 = $signed(wire359);
              reg364 <= (+(wire354[(1'h0):(1'h0)] ?
                  (!$unsigned(wire354[(1'h0):(1'h0)])) : reg363));
            end
          reg365 <= ($signed(((reg360 ?
                  $signed(reg361) : reg363) ^ (&{reg358}))) ?
              "GfMpxHd" : $signed("YXxXVpQ"));
        end
    end
  assign wire366 = $signed($signed({reg361[(2'h3):(1'h0)], "Qr"}));
  assign wire367 = reg364[(4'h8):(2'h3)];
  assign wire368 = wire357[(2'h2):(1'h0)];
  assign wire369 = reg362[(4'he):(4'hc)];
  assign wire370 = $unsigned($signed($signed((~&((8'hb5) ?
                       wire366 : reg365)))));
  assign wire371 = $unsigned(wire353);
  always
    @(posedge clk) begin
      for (forvar372 = (1'h0); (forvar372 < (2'h3)); forvar372 = (forvar372 + (1'h1)))
        begin
          if (((((wire370[(3'h4):(1'h0)] ?
                      (~&forvar372) : "64DfidaykSn9Zq4yOAJv7") ?
                  (wire356[(4'h8):(4'h8)] ?
                      $unsigned(wire369) : (wire356 ?
                          forvar372 : reg362)) : "NJ0ke15lOMGxnTnyeDPz") ?
              $unsigned((~|$signed(reg364))) : {$signed("AaCMW8nwQa09DHVskBwgMo")}) | $unsigned(wire359[(5'h14):(2'h2)])))
            begin
              reg373 = $unsigned($signed("IkzzcO2OJrRyq4vCFT"));
              reg374 <= $unsigned("neiumBvdmEcoq1oyMZM");
            end
          else
            begin
              reg373 <= ("Bxh6" <= $unsigned(reg364));
              reg374 <= (8'hb9);
              reg375 <= (|(($signed((~^wire354)) ^~ ($signed((8'hbd)) ?
                      (wire353 >>> (8'hb0)) : "uSygdx0v7eZpUSL0OXkBA")) ?
                  "KR59hrAF4SV0HoOP9rqEEk" : (&(^~(~&(8'h9f))))));
            end
        end
    end
  assign wire376 = "Xb";
  assign wire377 = $signed(reg361[(1'h1):(1'h0)]);
  assign wire378 = {"qapX"};
  assign wire379 = reg360;
  assign wire380 = wire370[(2'h3):(2'h3)];
  assign wire381 = (~&{$signed(forvar362[(2'h2):(1'h0)]), $unsigned(wire368)});
  assign wire382 = wire356;
  assign wire383 = $unsigned((!(($unsigned((7'h42)) & (reg358 ?
                       wire379 : reg360)) < $signed((~^wire353)))));
  assign wire384 = $unsigned({{"MAAsldGcPSLGBpekW", reg374}});
  assign wire385 = (+{wire381, "b8lXyuPgPGi2JdF"});
  assign wire386 = $unsigned($unsigned(reg358));
  always
    @(posedge clk) begin
      reg387 <= (~reg361);
      reg388 <= "8VXJ";
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module313  (y, clk, wire317, wire316, wire315, wire314);
  output wire [(32'h181):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'h9):(1'h0)] wire317;
  input wire signed [(4'hc):(1'h0)] wire316;
  input wire signed [(5'h14):(1'h0)] wire315;
  input wire signed [(4'hf):(1'h0)] wire314;
  reg [(4'hf):(1'h0)] reg348 = (1'h0);
  wire signed [(4'hd):(1'h0)] wire347;
  wire signed [(5'h10):(1'h0)] wire346;
  wire signed [(4'hf):(1'h0)] wire345;
  wire signed [(2'h3):(1'h0)] wire344;
  wire [(4'h9):(1'h0)] wire343;
  wire signed [(5'h16):(1'h0)] wire342;
  wire [(4'hb):(1'h0)] wire341;
  wire signed [(4'hb):(1'h0)] wire340;
  wire signed [(3'h7):(1'h0)] wire339;
  wire signed [(4'hd):(1'h0)] wire338;
  wire signed [(3'h5):(1'h0)] wire337;
  wire [(4'h8):(1'h0)] wire336;
  wire signed [(3'h7):(1'h0)] wire335;
  wire [(5'h16):(1'h0)] wire334;
  wire [(5'h16):(1'h0)] wire333;
  wire signed [(5'h13):(1'h0)] wire332;
  reg [(3'h4):(1'h0)] reg331 = (1'h0);
  reg signed [(4'he):(1'h0)] reg330 = (1'h0);
  reg [(4'h9):(1'h0)] reg329 = (1'h0);
  reg [(3'h5):(1'h0)] reg328 = (1'h0);
  reg [(4'hd):(1'h0)] reg327 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg326 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg325 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar324 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg322 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg321 = (1'h0);
  reg [(5'h15):(1'h0)] reg320 = (1'h0);
  reg [(5'h14):(1'h0)] reg319 = (1'h0);
  wire [(5'h16):(1'h0)] wire318;
  assign y = {reg348,
                 wire347,
                 wire346,
                 wire345,
                 wire344,
                 wire343,
                 wire342,
                 wire341,
                 wire340,
                 wire339,
                 wire338,
                 wire337,
                 wire336,
                 wire335,
                 wire334,
                 wire333,
                 wire332,
                 reg331,
                 reg330,
                 reg329,
                 reg328,
                 reg327,
                 reg326,
                 reg325,
                 forvar324,
                 reg323,
                 reg322,
                 reg321,
                 reg320,
                 reg319,
                 wire318,
                 (1'h0)};
  assign wire318 = "IfU1x1drawFmGn";
  always
    @(posedge clk) begin
      reg319 <= wire316[(2'h2):(1'h0)];
      if ($unsigned($signed($signed("1Nz1K4cyCQ"))))
        begin
          if ((("d1sCFv" ?
                  wire318[(2'h3):(2'h2)] : ((8'ha4) <= (^~(wire317 ~^ reg319)))) ?
              (7'h41) : "gyHAfybgQXr22UcC"))
            begin
              reg320 <= $signed((wire318[(5'h14):(3'h6)] ^ $unsigned(wire316)));
              reg321 = "Ci7iM";
            end
          else
            begin
              reg320 = ("FWa4qu" < wire317);
            end
          reg322 <= (~&wire318[(3'h5):(2'h3)]);
          reg323 <= reg321;
        end
      else
        begin
          reg320 <= ($unsigned((~{(reg322 ~^ reg323),
              (~wire314)})) ^ (~|(8'hbd)));
        end
      for (forvar324 = (1'h0); (forvar324 < (1'h1)); forvar324 = (forvar324 + (1'h1)))
        begin
          reg325 <= ((reg322 ?
              wire318[(3'h4):(1'h1)] : {($unsigned((8'hab)) - (!wire318)),
                  {(~&wire314)}}) <= "VT");
          if ("oiXqDGqKG")
            begin
              reg326 <= ($unsigned($unsigned($unsigned((reg322 >>> reg322)))) >>> (reg319[(4'hd):(2'h2)] ?
                  reg322 : ("r5d7grZuSRiNg" ?
                      ((^(8'hac)) ?
                          (reg325 ? wire314 : wire316) : ((8'ha1) ?
                              (8'hbe) : reg320)) : $signed((wire314 * wire315)))));
              reg327 <= $signed(reg325);
              reg328 <= reg323;
              reg329 = {"QuVkBd48x0dlrd44GfD", $signed($signed(reg327))};
            end
          else
            begin
              reg326 <= $signed(wire315);
              reg327 <= $signed("rIDkRHR0Cpi7S");
              reg328 <= {"vAUx31rDDV5TC"};
            end
        end
      reg330 <= $unsigned(reg329);
      reg331 <= {(^"4UwkIpMHz"), reg320[(3'h4):(3'h4)]};
    end
  assign wire332 = (~^wire318);
  assign wire333 = (reg321[(2'h2):(1'h0)] ?
                       $signed(reg320[(5'h14):(3'h4)]) : $unsigned((((~|(7'h44)) ?
                               {reg330} : ((7'h40) ? reg322 : (8'hac))) ?
                           reg328 : {$unsigned(reg327)})));
  assign wire334 = (8'ha5);
  assign wire335 = ((|reg331[(1'h0):(1'h0)]) >>> reg328[(1'h1):(1'h1)]);
  assign wire336 = ((^~(forvar324 ?
                       $unsigned("qzlqf") : ("TTXYla" ?
                           (wire334 ? (8'ha0) : wire335) : (reg329 ?
                               (7'h46) : reg322)))) | ((^~"BQgpXotOGnRHaBiHrA8t") ?
                       (~|"gn0N5Bg60sGJNnkW") : "uewiqPG2mS0maHd6A"));
  assign wire337 = $unsigned($signed($unsigned(($unsigned(reg326) <= "e2v5rFX64Ypx3k"))));
  assign wire338 = ("DO1LDp1" ? {(^forvar324[(1'h0):(1'h0)])} : "TY");
  assign wire339 = reg321[(4'hf):(3'h5)];
  assign wire340 = (|$unsigned({$unsigned({(8'hbb)}),
                       $signed($signed(reg321))}));
  assign wire341 = ((8'hb6) ?
                       $signed((wire335[(2'h3):(2'h3)] ?
                           ($unsigned(reg328) ?
                               "yskD2oBazA7xDK" : wire334) : $unsigned({reg321}))) : "tepHOwfAtAqO4BTwOz6");
  assign wire342 = ("p5Qe9RRwbc3" ?
                       (8'h9e) : (($unsigned($unsigned((8'hbc))) ?
                               (reg329[(2'h3):(2'h3)] ?
                                   ((8'hbe) + wire315) : (!(7'h40))) : reg327[(4'hc):(4'h8)]) ?
                           $unsigned((8'hae)) : $unsigned({$signed(reg330)})));
  assign wire343 = wire335[(1'h0):(1'h0)];
  assign wire344 = wire336;
  assign wire345 = ((reg322[(3'h4):(1'h1)] >= (^(^(8'hac)))) ?
                       "DpYusU9VFx" : "vi7oyJ1earcRL1CCb");
  assign wire346 = "rdOU5eSvJvQ6p7JGkq";
  assign wire347 = (7'h48);
  always
    @(posedge clk) begin
      reg348 <= $unsigned("a14woBJHseB");
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module200
#( parameter param247 = ((((((8'ha0) ? (7'h46) : (8'hac)) ? (~(8'hba)) : ((7'h46) ? (8'hb1) : (8'hb8))) >> (~(^(8'hb2)))) ? {(((8'ha6) < (8'hb1)) && ((7'h45) ? (8'hb4) : (7'h43))), (~((8'ha1) & (8'hb7)))} : (^~((^~(8'hac)) && {(8'h9e)}))) ? (((((8'hae) != (8'hb6)) ? (~(8'hb3)) : (~^(7'h40))) > ((^(7'h48)) ~^ ((8'ha4) > (8'hb5)))) << (((~&(8'hb8)) ? ((7'h42) ? (8'hbe) : (8'hb4)) : ((8'ha6) == (8'ha2))) ^~ (((8'ha0) ? (7'h40) : (8'ha8)) && (~|(8'h9c))))) : {{((^~(8'hb6)) ? (^~(8'hb9)) : ((8'ha6) ? (8'hae) : (8'hb2))), (-((8'hab) >>> (8'hab)))}})
, parameter param248 = param247 )
(y, clk, wire205, wire204, wire203, wire202, wire201);
  output wire [(32'h1e4):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire205;
  input wire [(5'h11):(1'h0)] wire204;
  input wire [(3'h6):(1'h0)] wire203;
  input wire [(5'h14):(1'h0)] wire202;
  input wire [(4'h8):(1'h0)] wire201;
  wire signed [(4'hf):(1'h0)] wire246;
  wire signed [(5'h16):(1'h0)] wire245;
  reg signed [(2'h3):(1'h0)] reg244 = (1'h0);
  wire signed [(4'h8):(1'h0)] wire243;
  wire [(3'h6):(1'h0)] wire242;
  wire signed [(4'hc):(1'h0)] wire241;
  wire signed [(5'h10):(1'h0)] wire240;
  reg [(4'h9):(1'h0)] reg239 = (1'h0);
  reg signed [(4'he):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar237 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg236 = (1'h0);
  reg [(5'h13):(1'h0)] reg235 = (1'h0);
  reg [(5'h17):(1'h0)] reg234 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg233 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg232 = (1'h0);
  reg [(4'hc):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg230 = (1'h0);
  reg [(4'hc):(1'h0)] reg229 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar228 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar227 = (1'h0);
  reg [(3'h6):(1'h0)] reg226 = (1'h0);
  reg [(4'he):(1'h0)] forvar225 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg224 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg223 = (1'h0);
  reg [(5'h12):(1'h0)] reg222 = (1'h0);
  reg [(5'h17):(1'h0)] reg221 = (1'h0);
  reg [(5'h14):(1'h0)] reg220 = (1'h0);
  reg [(3'h6):(1'h0)] reg219 = (1'h0);
  reg [(5'h12):(1'h0)] reg218 = (1'h0);
  reg [(3'h5):(1'h0)] forvar217 = (1'h0);
  reg [(3'h7):(1'h0)] forvar216 = (1'h0);
  wire signed [(4'hf):(1'h0)] wire215;
  wire signed [(3'h4):(1'h0)] wire214;
  wire [(5'h12):(1'h0)] wire213;
  wire signed [(5'h17):(1'h0)] wire212;
  wire signed [(3'h6):(1'h0)] wire211;
  wire signed [(3'h5):(1'h0)] wire210;
  wire [(4'h8):(1'h0)] wire209;
  wire [(3'h6):(1'h0)] wire208;
  wire signed [(3'h7):(1'h0)] wire207;
  wire [(4'hf):(1'h0)] wire206;
  assign y = {wire246,
                 wire245,
                 reg244,
                 wire243,
                 wire242,
                 wire241,
                 wire240,
                 reg239,
                 reg238,
                 forvar237,
                 reg236,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg230,
                 reg229,
                 forvar228,
                 forvar227,
                 reg226,
                 forvar225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg219,
                 reg218,
                 forvar217,
                 forvar216,
                 wire215,
                 wire214,
                 wire213,
                 wire212,
                 wire211,
                 wire210,
                 wire209,
                 wire208,
                 wire207,
                 wire206,
                 (1'h0)};
  assign wire206 = wire204[(4'h8):(1'h1)];
  assign wire207 = ($signed(wire205[(2'h3):(2'h2)]) > wire204[(3'h7):(3'h5)]);
  assign wire208 = {(|"xnC2NK4")};
  assign wire209 = (~wire203[(3'h5):(3'h4)]);
  assign wire210 = $unsigned({$signed(((wire209 * wire209) ?
                           wire201 : wire205)),
                       ((wire201[(3'h6):(1'h1)] ?
                           $signed((8'ha8)) : "VME7CgsPfk4") < (&$signed(wire205)))});
  assign wire211 = (8'hbb);
  assign wire212 = "JtB";
  assign wire213 = (($signed(wire204) ? (8'hba) : wire211) ?
                       ("2tv0rbYPlXWg5mbG5J" >> wire209) : $signed("XPsQCClbni4"));
  assign wire214 = ({(8'hb5),
                       $signed($unsigned(wire207[(3'h7):(3'h5)]))} >= $signed($unsigned((~|((8'hbf) ?
                       wire204 : wire208)))));
  assign wire215 = $unsigned((^~$unsigned($signed({wire213, (8'hb6)}))));
  always
    @(posedge clk) begin
      for (forvar216 = (1'h0); (forvar216 < (3'h4)); forvar216 = (forvar216 + (1'h1)))
        begin
          for (forvar217 = (1'h0); (forvar217 < (2'h3)); forvar217 = (forvar217 + (1'h1)))
            begin
              reg218 <= wire202[(4'he):(2'h2)];
              reg219 <= (wire207[(1'h0):(1'h0)] ?
                  {"ZLSt1MALBDD1vKwaara",
                      wire202} : (~$unsigned(wire209[(3'h5):(1'h1)])));
              reg220 <= $signed(wire215[(4'he):(1'h0)]);
              reg221 <= (7'h44);
            end
          reg222 <= $signed((^~(^~$signed((7'h43)))));
          reg223 = $signed("9WQ7l7fOMXdkfnh3Fze5");
          reg224 <= reg220[(1'h0):(1'h0)];
          for (forvar225 = (1'h0); (forvar225 < (3'h4)); forvar225 = (forvar225 + (1'h1)))
            begin
              reg226 <= $signed(wire210[(2'h3):(1'h0)]);
            end
        end
      for (forvar227 = (1'h0); (forvar227 < (3'h4)); forvar227 = (forvar227 + (1'h1)))
        begin
          for (forvar228 = (1'h0); (forvar228 < (1'h1)); forvar228 = (forvar228 + (1'h1)))
            begin
              reg229 <= wire214;
              reg230 <= wire211;
              reg231 = $signed(forvar228[(2'h2):(1'h1)]);
              reg232 <= reg218[(3'h6):(1'h1)];
            end
          reg233 <= $unsigned(((((8'hba) ?
                  reg219[(3'h4):(3'h4)] : forvar217[(1'h0):(1'h0)]) & (8'hb4)) ?
              (reg231 == "k07l7sgc") : "y"));
          reg234 <= "mJkWn21bCJQ93FOUCu";
        end
      reg235 <= (wire215[(3'h4):(2'h2)] ? (~&reg220) : reg233[(1'h1):(1'h1)]);
      reg236 <= (&(^(reg222[(3'h4):(1'h0)] ?
          reg220[(4'he):(3'h4)] : $signed((reg230 ? wire209 : (8'ha3))))));
      for (forvar237 = (1'h0); (forvar237 < (2'h3)); forvar237 = (forvar237 + (1'h1)))
        begin
          reg238 = $signed(reg226);
          reg239 = {reg233[(3'h5):(1'h1)],
              $signed(($signed("FeVENI1") ?
                  reg230 : (+forvar227[(3'h7):(2'h2)])))};
        end
    end
  assign wire240 = wire201[(1'h0):(1'h0)];
  assign wire241 = wire211;
  assign wire242 = {("BW9" ?
                           ($signed({wire215}) ?
                               $unsigned($unsigned(reg219)) : $signed((~^reg226))) : wire210[(1'h0):(1'h0)])};
  assign wire243 = (^{(-(~^$unsigned(wire207)))});
  always
    @(posedge clk) begin
      reg244 <= (((~reg231) + ($unsigned($signed(wire208)) <<< ((reg224 ^~ reg236) >= (reg234 + reg236)))) ?
          "D5dpKRG" : $unsigned(wire203));
    end
  assign wire245 = $signed((reg220 - (forvar225[(1'h0):(1'h0)] ?
                       (wire207[(3'h4):(2'h2)] ?
                           forvar228 : (reg233 == reg226)) : ((~|reg235) ?
                           $unsigned(reg219) : (~&reg219)))));
  assign wire246 = (~^$signed($unsigned({$signed(wire207)})));
endmodule