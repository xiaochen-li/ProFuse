(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param710 = {{(((^~(8'hba)) <<< (^~(8'h9d))) ? {((8'ha7) ? (8'hb6) : (8'haa)), ((8'haa) ? (8'hb1) : (8'hb8))} : ((+(8'ha1)) ? (~&(7'h42)) : ((8'hb6) ? (8'hb3) : (8'ha1))))}, ((((~(8'hba)) && {(7'h44), (7'h42)}) <<< {((8'hba) <= (8'ha1)), ((8'hba) ? (8'hba) : (7'h41))}) ? ((|(~(8'hb8))) ? (((8'hb6) == (8'hb8)) ? ((8'haa) ? (7'h44) : (8'hb0)) : {(8'haf)}) : ((-(8'ha1)) ? ((8'hbd) ? (8'hb7) : (8'hb2)) : ((8'haa) && (8'hb3)))) : (^~((~^(8'had)) && ((7'h40) == (7'h44)))))})
(y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h3ed):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire0;
  input wire signed [(3'h4):(1'h0)] wire1;
  input wire signed [(4'h9):(1'h0)] wire2;
  input wire [(5'h10):(1'h0)] wire3;
  wire [(5'h13):(1'h0)] wire709;
  wire [(3'h5):(1'h0)] wire687;
  wire signed [(2'h2):(1'h0)] wire685;
  wire signed [(2'h3):(1'h0)] wire684;
  wire signed [(5'h13):(1'h0)] wire683;
  wire signed [(4'he):(1'h0)] wire679;
  wire [(3'h7):(1'h0)] wire678;
  wire [(5'h11):(1'h0)] wire641;
  wire [(4'hd):(1'h0)] wire4;
  wire signed [(4'hf):(1'h0)] wire5;
  wire signed [(4'h9):(1'h0)] wire15;
  wire signed [(3'h5):(1'h0)] wire639;
  wire signed [(2'h3):(1'h0)] wire674;
  wire signed [(4'h9):(1'h0)] wire675;
  wire [(3'h7):(1'h0)] wire676;
  wire signed [(3'h5):(1'h0)] wire681;
  wire signed [(5'h12):(1'h0)] wire689;
  wire [(5'h12):(1'h0)] wire707;
  reg [(3'h5):(1'h0)] reg704 = (1'h0);
  reg [(2'h3):(1'h0)] reg702 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg701 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg700 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg697 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg696 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg691 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg672 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg670 = (1'h0);
  reg [(4'ha):(1'h0)] reg669 = (1'h0);
  reg [(5'h10):(1'h0)] reg668 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg667 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg665 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg659 = (1'h0);
  reg [(4'hf):(1'h0)] reg658 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg654 = (1'h0);
  reg [(4'hc):(1'h0)] reg651 = (1'h0);
  reg [(5'h13):(1'h0)] reg648 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg646 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg9 = (1'h0);
  reg [(3'h4):(1'h0)] reg10 = (1'h0);
  reg [(5'h10):(1'h0)] reg11 = (1'h0);
  reg [(4'he):(1'h0)] reg13 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg16 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg19 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg20 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg21 = (1'h0);
  reg [(5'h12):(1'h0)] reg24 = (1'h0);
  reg [(5'h13):(1'h0)] reg25 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg26 = (1'h0);
  reg [(4'hc):(1'h0)] reg706 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg705 = (1'h0);
  reg [(3'h6):(1'h0)] forvar703 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg699 = (1'h0);
  reg [(4'hd):(1'h0)] forvar698 = (1'h0);
  reg [(3'h6):(1'h0)] forvar695 = (1'h0);
  reg [(5'h10):(1'h0)] reg694 = (1'h0);
  reg [(4'hb):(1'h0)] reg693 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar692 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar690 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg686 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg673 = (1'h0);
  reg [(3'h7):(1'h0)] reg671 = (1'h0);
  reg [(4'hd):(1'h0)] forvar666 = (1'h0);
  reg [(4'hd):(1'h0)] reg664 = (1'h0);
  reg [(5'h11):(1'h0)] reg663 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg662 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg661 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar660 = (1'h0);
  reg [(3'h7):(1'h0)] reg657 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar656 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar655 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg653 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg652 = (1'h0);
  reg [(4'hf):(1'h0)] reg650 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar649 = (1'h0);
  reg [(4'hb):(1'h0)] reg647 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg645 = (1'h0);
  reg [(5'h12):(1'h0)] forvar644 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar643 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg22 = (1'h0);
  reg [(5'h15):(1'h0)] forvar18 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg17 = (1'h0);
  reg [(3'h4):(1'h0)] reg14 = (1'h0);
  reg [(5'h11):(1'h0)] reg12 = (1'h0);
  reg [(4'h8):(1'h0)] reg8 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar7 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar6 = (1'h0);
  assign y = {wire709,
                 wire687,
                 wire685,
                 wire684,
                 wire683,
                 wire679,
                 wire678,
                 wire641,
                 wire4,
                 wire5,
                 wire15,
                 wire639,
                 wire674,
                 wire675,
                 wire676,
                 wire681,
                 wire689,
                 wire707,
                 reg704,
                 reg702,
                 reg701,
                 reg700,
                 reg697,
                 reg696,
                 reg691,
                 reg672,
                 reg670,
                 reg669,
                 reg668,
                 reg667,
                 reg665,
                 reg659,
                 reg658,
                 reg654,
                 reg651,
                 reg648,
                 reg646,
                 reg9,
                 reg10,
                 reg11,
                 reg13,
                 reg16,
                 reg19,
                 reg20,
                 reg21,
                 reg24,
                 reg25,
                 reg26,
                 reg706,
                 reg705,
                 forvar703,
                 reg699,
                 forvar698,
                 forvar695,
                 reg694,
                 reg693,
                 forvar692,
                 forvar690,
                 reg686,
                 reg673,
                 reg671,
                 forvar666,
                 reg664,
                 reg663,
                 reg662,
                 reg661,
                 forvar660,
                 reg657,
                 forvar656,
                 forvar655,
                 reg653,
                 reg652,
                 reg650,
                 forvar649,
                 reg647,
                 reg645,
                 forvar644,
                 forvar643,
                 reg23,
                 reg22,
                 forvar18,
                 reg17,
                 reg14,
                 reg12,
                 reg8,
                 forvar7,
                 forvar6,
                 (1'h0)};
  assign wire4 = wire2;
  assign wire5 = wire2;
  always
    @(posedge clk) begin
      for (forvar6 = (1'h0); (forvar6 < (1'h0)); forvar6 = (forvar6 + (1'h1)))
        begin
          for (forvar7 = (1'h0); (forvar7 < (3'h4)); forvar7 = (forvar7 + (1'h1)))
            begin
              reg8 = forvar7;
              reg9 <= wire0[(2'h3):(2'h3)];
              reg10 <= {((+reg9[(4'hf):(4'h8)]) ?
                      (((~reg8) != (wire0 * forvar7)) ?
                          (wire0[(1'h1):(1'h0)] <= (~^reg9)) : wire2[(2'h3):(1'h0)]) : (wire2 <<< ($signed(wire3) ~^ $signed(reg9))))};
              reg11 <= $signed($unsigned(wire1[(2'h2):(2'h2)]));
            end
        end
      reg12 = wire3[(2'h3):(2'h3)];
      reg13 <= ((&$unsigned("K2oaJmhS8K71BMvsD2")) ?
          reg11 : (&wire5[(3'h4):(2'h2)]));
      reg14 = (8'hb6);
    end
  assign wire15 = $signed(wire2);
  always
    @(posedge clk) begin
      reg16 <= reg13[(4'h8):(3'h6)];
      reg17 = (wire15[(2'h2):(2'h2)] <= (reg9 <= (^~wire0)));
      for (forvar18 = (1'h0); (forvar18 < (3'h4)); forvar18 = (forvar18 + (1'h1)))
        begin
          reg19 <= $signed($unsigned((&reg17[(4'h8):(2'h2)])));
          reg20 <= (((8'hb7) && (($unsigned((8'hb9)) ?
                  "u2ExMpnUVcywf0Q" : (-forvar18)) || $unsigned($signed(wire2)))) ?
              (wire5 >> wire15) : "RVsbFpeqO9m");
          if ((reg16[(3'h4):(1'h0)] ?
              ((7'h41) ?
                  {$signed($unsigned(reg20))} : wire0[(5'h14):(2'h2)]) : ((~((8'hbf) < $unsigned(wire15))) ?
                  (reg11[(2'h3):(2'h2)] & ($signed(wire4) >= (reg11 ?
                      (7'h44) : (8'hb2)))) : $signed(reg16))))
            begin
              reg21 <= forvar18;
              reg22 = $signed($unsigned({((8'had) ?
                      {wire5} : $unsigned(reg10))}));
              reg23 = wire15[(3'h4):(2'h3)];
            end
          else
            begin
              reg21 <= reg11;
              reg24 <= $unsigned(reg9);
              reg25 <= (^~((("DBnqWy5Y4cTse" == $signed(reg11)) ?
                  reg24[(2'h3):(1'h0)] : (wire5 >= $unsigned(reg23))) || wire5[(3'h7):(3'h7)]));
            end
        end
      reg26 <= reg19;
    end
  module27 #() modinst640 (.wire31(reg11), .wire32(wire0), .clk(clk), .wire28(reg25), .wire29(reg16), .y(wire639), .wire30(reg9));
  module477 #() modinst642 (.y(wire641), .wire480(reg25), .wire479(reg24), .wire481(reg20), .wire478(wire2), .clk(clk));
  always
    @(posedge clk) begin
      for (forvar643 = (1'h0); (forvar643 < (2'h2)); forvar643 = (forvar643 + (1'h1)))
        begin
          for (forvar644 = (1'h0); (forvar644 < (1'h1)); forvar644 = (forvar644 + (1'h1)))
            begin
              reg645 = ($unsigned(forvar643[(3'h6):(2'h3)]) != (wire3[(1'h1):(1'h1)] ?
                  $unsigned(($unsigned(reg11) ?
                      reg10[(2'h2):(1'h0)] : ((8'hac) ?
                          reg26 : wire4))) : reg24));
              reg646 <= $signed(reg11[(4'hf):(4'hb)]);
              reg647 = (^wire641);
              reg648 <= reg21;
            end
          for (forvar649 = (1'h0); (forvar649 < (1'h1)); forvar649 = (forvar649 + (1'h1)))
            begin
              reg650 = {(reg21[(3'h7):(3'h7)] ?
                      forvar649[(1'h0):(1'h0)] : reg21)};
              reg651 <= reg16;
              reg652 = {$unsigned({((&reg645) + reg650),
                      (|reg648[(1'h1):(1'h0)])}),
                  reg645[(1'h1):(1'h1)]};
              reg653 = reg24[(3'h6):(3'h4)];
              reg654 <= {$signed("3d6CcI"),
                  (((+"bpl9XlGMsi") >>> (~(forvar643 << wire4))) & reg10)};
            end
        end
      for (forvar655 = (1'h0); (forvar655 < (1'h1)); forvar655 = (forvar655 + (1'h1)))
        begin
          for (forvar656 = (1'h0); (forvar656 < (2'h3)); forvar656 = (forvar656 + (1'h1)))
            begin
              reg657 = (forvar644[(3'h6):(1'h0)] & reg645[(4'hd):(2'h3)]);
            end
          reg658 <= (|"t");
          reg659 <= (^~(~&{(wire3[(1'h1):(1'h0)] >= (reg10 * (8'hae))),
              (+$unsigned(reg651))}));
        end
      for (forvar660 = (1'h0); (forvar660 < (1'h0)); forvar660 = (forvar660 + (1'h1)))
        begin
          if (({$signed($unsigned((reg21 ? (8'h9d) : reg650))),
                  ($unsigned("HpHMGX2JJAawU") > $signed((reg652 ?
                      reg20 : reg659)))} ?
              forvar655 : forvar655))
            begin
              reg661 = $signed(wire4);
              reg662 = forvar660[(2'h3):(2'h2)];
              reg663 = forvar655[(4'hc):(1'h0)];
              reg664 = reg657;
              reg665 <= (&$unsigned($signed(reg653)));
            end
          else
            begin
              reg661 = ($unsigned(wire0[(5'h11):(4'h9)]) ?
                  reg659 : $signed((~&wire4[(2'h3):(1'h0)])));
            end
          for (forvar666 = (1'h0); (forvar666 < (1'h0)); forvar666 = (forvar666 + (1'h1)))
            begin
              reg667 <= reg647[(4'h9):(3'h7)];
              reg668 <= $signed(reg665);
              reg669 <= (~|(forvar655[(3'h7):(1'h1)] ^~ reg26));
              reg670 <= $unsigned((!reg662[(3'h6):(3'h5)]));
              reg671 = ((({(~&forvar655)} ?
                      {wire639[(1'h0):(1'h0)],
                          $unsigned((8'hbd))} : (^(|reg16))) ?
                  ($unsigned((reg668 ?
                      reg653 : wire2)) ~^ $unsigned($unsigned(wire2))) : (8'hb5)) && ((^reg653[(4'hd):(3'h4)]) ?
                  reg20 : (~reg21)));
            end
          reg672 <= reg648[(2'h3):(2'h2)];
        end
      reg673 = reg659;
    end
  assign wire674 = reg654;
  assign wire675 = wire0[(5'h10):(3'h4)];
  module27 #() modinst677 (wire676, clk, reg25, wire3, reg668, reg9, reg20);
  assign wire678 = $unsigned((((8'ha1) <<< ((^reg13) * $signed((8'hb3)))) << (reg20 ?
                       "3NLBITVM0" : (wire2 ? (wire0 == reg651) : (!wire0)))));
  module65 #() modinst680 (wire679, clk, reg11, reg669, reg648, reg668, wire0);
  module65 #() modinst682 (wire681, clk, reg21, reg648, reg16, wire675, reg659);
  assign wire683 = ((((8'ha7) ?
                           wire674[(2'h2):(2'h2)] : $signed(wire681)) + reg659[(5'h13):(5'h11)]) ?
                       $unsigned(reg667[(2'h3):(1'h1)]) : reg659);
  assign wire684 = reg648[(4'hd):(4'h8)];
  assign wire685 = (((reg26[(4'h9):(3'h6)] ? (^(~(8'h9f))) : wire676) ?
                       ($unsigned((~|reg16)) ?
                           (!reg654[(1'h1):(1'h1)]) : (reg648 * (reg20 ?
                               wire15 : wire676))) : (($signed(wire683) >>> wire681[(3'h4):(3'h4)]) <= (~wire676[(3'h5):(2'h3)]))) > {((((8'hb9) + (8'hb0)) ?
                               (^reg651) : wire679[(1'h1):(1'h1)]) ?
                           reg658[(2'h3):(1'h1)] : ((reg648 + wire1) != (&(8'hbe))))});
  always
    @(posedge clk) begin
      reg686 = {reg24[(4'ha):(1'h1)]};
    end
  module65 #() modinst688 (.wire68(reg658), .wire66(reg648), .wire67(wire641), .wire70(reg669), .wire69(reg9), .y(wire687), .clk(clk));
  assign wire689 = ({($signed($unsigned(wire15)) ^ $signed($signed(reg19)))} ^ (($signed($signed(reg20)) ~^ ($unsigned(reg651) ?
                           wire15 : (wire3 <<< reg648))) ?
                       $unsigned("Caz2DLFBkXXGK9") : $signed(wire687[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      for (forvar690 = (1'h0); (forvar690 < (2'h3)); forvar690 = (forvar690 + (1'h1)))
        begin
          reg691 <= reg669[(3'h7):(3'h4)];
          for (forvar692 = (1'h0); (forvar692 < (2'h3)); forvar692 = (forvar692 + (1'h1)))
            begin
              reg693 = reg20[(2'h2):(1'h0)];
              reg694 = {({$signed($unsigned(wire683)),
                          $signed((reg26 ? reg21 : reg651))} ?
                      (!$unsigned($signed(reg648))) : ((~^$unsigned(reg13)) ?
                          (|(+reg25)) : wire5)),
                  reg16[(5'h11):(4'hb)]};
            end
          for (forvar695 = (1'h0); (forvar695 < (3'h4)); forvar695 = (forvar695 + (1'h1)))
            begin
              reg696 <= (~^wire676);
              reg697 <= $signed({$signed((~$unsigned(reg21))),
                  $unsigned($unsigned({wire5}))});
            end
          for (forvar698 = (1'h0); (forvar698 < (1'h0)); forvar698 = (forvar698 + (1'h1)))
            begin
              reg699 = {wire3[(4'hb):(3'h7)]};
              reg700 <= $signed(reg691[(3'h4):(2'h3)]);
              reg701 <= (|($signed({reg693[(4'h8):(3'h4)],
                  (-reg699)}) & $signed(reg669)));
            end
          reg702 <= {$signed(({(forvar692 >>> (8'hb7)),
                  (reg19 == (8'hb3))} && reg26))};
        end
      for (forvar703 = (1'h0); (forvar703 < (2'h2)); forvar703 = (forvar703 + (1'h1)))
        begin
          reg704 <= (^~$signed((wire2 ?
              (8'hbe) : (reg648 ? wire689 : wire676[(2'h2):(2'h2)]))));
        end
      reg705 = {{(8'ha9)},
          $unsigned((reg11[(3'h4):(3'h4)] + reg646[(2'h3):(2'h3)]))};
      reg706 = reg21[(1'h1):(1'h0)];
    end
  module65 #() modinst708 (.wire69(reg19), .clk(clk), .wire66(wire683), .wire70(reg672), .wire68(wire0), .y(wire707), .wire67(wire5));
  assign wire709 = reg659[(2'h3):(2'h3)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module27
#(parameter param638 = ((((((8'hb6) ? (7'h44) : (8'hbf)) > {(8'ha3), (8'hbd)}) ? ((~|(8'hb4)) ^ ((8'ha7) - (8'ha1))) : (^((8'hab) ? (8'hac) : (8'ha2)))) ? (^~((~^(8'hbe)) ? (^(8'ha8)) : (~|(8'hb2)))) : ((((8'h9f) == (8'hbb)) & (~&(8'hb1))) ? ((^~(8'hb5)) ? {(8'ha5), (8'hb2)} : ((8'ha3) ? (8'ha9) : (8'hb2))) : ((-(8'hbb)) ? ((8'hbe) ? (8'hb3) : (8'ha1)) : ((8'h9c) == (7'h44))))) == (({((8'hbf) ? (8'ha2) : (8'ha8))} <= ((!(8'hbc)) * {(7'h43)})) == ((8'ha2) ? (((8'hab) ? (7'h41) : (8'ha1)) ? ((8'ha7) ? (8'hbf) : (8'hb8)) : (~^(8'hac))) : (((8'h9c) && (8'ha2)) <= {(8'hbf), (8'hb6)})))))
(y, clk, wire32, wire31, wire30, wire29, wire28);
  output wire [(32'h5ef):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire32;
  input wire signed [(5'h10):(1'h0)] wire31;
  input wire [(5'h10):(1'h0)] wire30;
  input wire signed [(4'h9):(1'h0)] wire29;
  input wire [(5'h13):(1'h0)] wire28;
  wire [(5'h14):(1'h0)] wire385;
  wire [(5'h11):(1'h0)] wire273;
  wire [(4'ha):(1'h0)] wire171;
  wire [(5'h14):(1'h0)] wire170;
  wire [(4'hd):(1'h0)] wire169;
  wire [(4'ha):(1'h0)] wire167;
  wire signed [(4'hf):(1'h0)] wire407;
  wire [(4'hf):(1'h0)] wire408;
  wire [(5'h14):(1'h0)] wire471;
  wire [(4'he):(1'h0)] wire473;
  wire signed [(3'h7):(1'h0)] wire474;
  wire signed [(4'he):(1'h0)] wire475;
  wire signed [(3'h5):(1'h0)] wire476;
  wire signed [(4'hc):(1'h0)] wire583;
  reg [(4'hc):(1'h0)] reg637 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg636 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg635 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg634 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg629 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg627 = (1'h0);
  reg [(4'hd):(1'h0)] reg626 = (1'h0);
  reg [(4'hc):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg617 = (1'h0);
  reg [(5'h12):(1'h0)] reg616 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg613 = (1'h0);
  reg [(3'h7):(1'h0)] reg612 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg608 = (1'h0);
  reg [(4'h8):(1'h0)] reg607 = (1'h0);
  reg [(4'hb):(1'h0)] reg605 = (1'h0);
  reg [(3'h6):(1'h0)] reg604 = (1'h0);
  reg [(5'h11):(1'h0)] reg602 = (1'h0);
  reg signed [(4'he):(1'h0)] reg600 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg596 = (1'h0);
  reg [(4'h9):(1'h0)] reg595 = (1'h0);
  reg [(4'h8):(1'h0)] reg593 = (1'h0);
  reg [(3'h6):(1'h0)] reg592 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg591 = (1'h0);
  reg [(3'h6):(1'h0)] reg405 = (1'h0);
  reg [(5'h15):(1'h0)] reg402 = (1'h0);
  reg [(5'h12):(1'h0)] reg401 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg400 = (1'h0);
  reg [(5'h11):(1'h0)] reg399 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg390 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg395 = (1'h0);
  reg [(3'h6):(1'h0)] reg393 = (1'h0);
  reg [(5'h14):(1'h0)] reg387 = (1'h0);
  reg [(4'hc):(1'h0)] reg35 = (1'h0);
  reg [(4'hc):(1'h0)] reg37 = (1'h0);
  reg [(5'h10):(1'h0)] reg39 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg45 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg47 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg48 = (1'h0);
  reg [(4'hb):(1'h0)] reg49 = (1'h0);
  reg [(4'hf):(1'h0)] reg52 = (1'h0);
  reg [(5'h15):(1'h0)] reg53 = (1'h0);
  reg [(4'hf):(1'h0)] reg55 = (1'h0);
  reg [(5'h15):(1'h0)] reg56 = (1'h0);
  reg [(4'hc):(1'h0)] reg57 = (1'h0);
  reg [(4'ha):(1'h0)] reg58 = (1'h0);
  reg [(5'h15):(1'h0)] reg62 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg63 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg51 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg633 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg632 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg631 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg630 = (1'h0);
  reg signed [(4'he):(1'h0)] reg628 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg623 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg622 = (1'h0);
  reg [(4'hb):(1'h0)] reg621 = (1'h0);
  reg [(4'hf):(1'h0)] reg620 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar619 = (1'h0);
  reg [(4'h8):(1'h0)] forvar618 = (1'h0);
  reg [(5'h15):(1'h0)] reg615 = (1'h0);
  reg [(4'ha):(1'h0)] forvar614 = (1'h0);
  reg [(4'hd):(1'h0)] reg611 = (1'h0);
  reg [(3'h4):(1'h0)] reg610 = (1'h0);
  reg [(3'h6):(1'h0)] reg609 = (1'h0);
  reg [(5'h14):(1'h0)] reg606 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar606 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg603 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg601 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg599 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg598 = (1'h0);
  reg [(4'he):(1'h0)] forvar597 = (1'h0);
  reg [(5'h10):(1'h0)] reg594 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg590 = (1'h0);
  reg [(5'h13):(1'h0)] reg589 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar588 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg587 = (1'h0);
  reg [(2'h2):(1'h0)] forvar586 = (1'h0);
  reg [(4'hf):(1'h0)] forvar585 = (1'h0);
  reg [(4'hd):(1'h0)] reg406 = (1'h0);
  reg [(5'h15):(1'h0)] forvar404 = (1'h0);
  reg [(4'hb):(1'h0)] forvar403 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg398 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar397 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar392 = (1'h0);
  reg [(4'hb):(1'h0)] forvar387 = (1'h0);
  reg [(3'h4):(1'h0)] reg396 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg394 = (1'h0);
  reg [(3'h6):(1'h0)] reg392 = (1'h0);
  reg [(4'hd):(1'h0)] reg391 = (1'h0);
  reg [(4'h8):(1'h0)] forvar390 = (1'h0);
  reg [(3'h4):(1'h0)] reg389 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg388 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg54 = (1'h0);
  reg [(2'h2):(1'h0)] forvar52 = (1'h0);
  reg [(5'h10):(1'h0)] reg46 = (1'h0);
  reg [(5'h10):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg61 = (1'h0);
  reg [(3'h5):(1'h0)] reg60 = (1'h0);
  reg [(5'h10):(1'h0)] reg59 = (1'h0);
  reg [(4'hc):(1'h0)] forvar54 = (1'h0);
  reg [(3'h5):(1'h0)] forvar51 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg50 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar46 = (1'h0);
  reg [(4'hb):(1'h0)] reg44 = (1'h0);
  reg [(5'h10):(1'h0)] reg43 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg41 = (1'h0);
  reg [(5'h11):(1'h0)] reg40 = (1'h0);
  reg [(3'h6):(1'h0)] reg38 = (1'h0);
  reg [(3'h4):(1'h0)] forvar36 = (1'h0);
  reg [(5'h14):(1'h0)] reg34 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg33 = (1'h0);
  assign y = {wire385,
                 wire273,
                 wire171,
                 wire170,
                 wire169,
                 wire167,
                 wire407,
                 wire408,
                 wire471,
                 wire473,
                 wire474,
                 wire475,
                 wire476,
                 wire583,
                 reg637,
                 reg636,
                 reg635,
                 reg634,
                 reg629,
                 reg627,
                 reg626,
                 reg625,
                 reg617,
                 reg616,
                 reg613,
                 reg612,
                 reg608,
                 reg607,
                 reg605,
                 reg604,
                 reg602,
                 reg600,
                 reg596,
                 reg595,
                 reg593,
                 reg592,
                 reg591,
                 reg405,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg390,
                 reg395,
                 reg393,
                 reg387,
                 reg35,
                 reg37,
                 reg39,
                 reg45,
                 reg47,
                 reg48,
                 reg49,
                 reg52,
                 reg53,
                 reg55,
                 reg56,
                 reg57,
                 reg58,
                 reg62,
                 reg63,
                 reg51,
                 reg633,
                 reg632,
                 reg631,
                 reg630,
                 reg628,
                 reg624,
                 reg623,
                 reg622,
                 reg621,
                 reg620,
                 forvar619,
                 forvar618,
                 reg615,
                 forvar614,
                 reg611,
                 reg610,
                 reg609,
                 reg606,
                 forvar606,
                 reg603,
                 reg601,
                 reg599,
                 reg598,
                 forvar597,
                 reg594,
                 reg590,
                 reg589,
                 forvar588,
                 reg587,
                 forvar586,
                 forvar585,
                 reg406,
                 forvar404,
                 forvar403,
                 reg398,
                 forvar397,
                 forvar392,
                 forvar387,
                 reg396,
                 reg394,
                 reg392,
                 reg391,
                 forvar390,
                 reg389,
                 reg388,
                 reg54,
                 forvar52,
                 reg46,
                 reg64,
                 reg61,
                 reg60,
                 reg59,
                 forvar54,
                 forvar51,
                 reg50,
                 forvar46,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg38,
                 forvar36,
                 reg34,
                 reg33,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg33 = wire31[(4'hd):(2'h2)];
    end
  always
    @(posedge clk) begin
      reg34 = {$signed(wire32[(3'h7):(3'h5)]),
          (^(((8'h9e) ? (wire31 ? wire30 : (8'hb1)) : {wire31}) ?
              $unsigned(((8'had) < wire30)) : (-(wire32 | wire28))))};
      reg35 <= wire32[(3'h7):(3'h4)];
      for (forvar36 = (1'h0); (forvar36 < (2'h2)); forvar36 = (forvar36 + (1'h1)))
        begin
          reg37 <= wire32;
          if (reg37[(3'h6):(3'h6)])
            begin
              reg38 = $signed(reg34[(4'h9):(3'h4)]);
              reg39 <= $unsigned({$signed((~^reg37[(1'h0):(1'h0)]))});
              reg40 = (-(wire29 + reg35));
              reg41 = {$unsigned((^~($unsigned(forvar36) & $signed(forvar36))))};
              reg42 = (wire30[(3'h4):(2'h3)] == "DgO2ER139Tk3");
            end
          else
            begin
              reg38 = ($signed({reg37}) | $signed((((reg40 ?
                  wire28 : wire30) ^~ (~&reg37)) != ({reg37} ?
                  (reg41 ? wire31 : reg41) : (8'ha1)))));
              reg40 = wire32[(3'h4):(2'h3)];
            end
          reg43 = $unsigned($unsigned((8'hae)));
          reg44 = $signed((reg42[(2'h3):(1'h0)] * ($signed((wire29 ?
              (8'haa) : reg40)) ^ $signed($unsigned(wire29)))));
        end
      reg45 <= $unsigned(($unsigned("tRLNxqlK18O") ?
          $unsigned($signed($unsigned(wire28))) : $unsigned(((&reg41) ?
              $signed(reg42) : $signed(forvar36)))));
      if ((&reg42))
        begin
          for (forvar46 = (1'h0); (forvar46 < (1'h1)); forvar46 = (forvar46 + (1'h1)))
            begin
              reg47 <= $unsigned(reg42);
              reg48 <= reg45;
              reg49 <= reg48;
              reg50 = {reg43};
            end
          for (forvar51 = (1'h0); (forvar51 < (1'h1)); forvar51 = (forvar51 + (1'h1)))
            begin
              reg52 <= reg41[(2'h2):(1'h1)];
              reg53 <= wire31[(3'h5):(1'h1)];
            end
          for (forvar54 = (1'h0); (forvar54 < (1'h0)); forvar54 = (forvar54 + (1'h1)))
            begin
              reg55 <= "Jie0U";
              reg56 <= reg53;
              reg57 <= $signed($signed($signed(reg52[(4'hb):(3'h6)])));
              reg58 <= ((reg38 & (~&"pY")) ?
                  wire31 : $unsigned((reg38 ?
                      reg56[(5'h13):(4'hf)] : (-reg55[(2'h3):(2'h3)]))));
            end
          reg59 = (~|$signed((+$signed({reg44}))));
          if ((+$unsigned((^(+$unsigned(reg42))))))
            begin
              reg60 = wire32[(2'h3):(2'h2)];
              reg61 = ($signed($unsigned($signed((~reg56)))) ?
                  (wire32[(2'h3):(2'h2)] ?
                      (wire28 ?
                          ((^forvar46) != reg40[(4'h9):(3'h4)]) : ((reg40 * reg52) ?
                              reg43 : reg34[(3'h7):(3'h6)])) : (({reg58,
                              reg39} - reg45) ?
                          forvar36 : ($signed(wire31) << (reg56 ?
                              forvar51 : reg41)))) : ("nVugZFIgquW" && (((reg53 ?
                          reg58 : reg59) && reg47[(1'h1):(1'h0)]) ?
                      $unsigned((~|(8'hbb))) : reg35)));
            end
          else
            begin
              reg62 <= (^(reg56[(5'h15):(3'h5)] | {$signed($unsigned(wire28)),
                  (-reg45[(2'h2):(2'h2)])}));
              reg63 <= $signed("prGiaU19POee8m");
              reg64 = ($unsigned((((^reg57) == (^~reg60)) || (reg49 ?
                  reg61 : (8'ha6)))) >= $unsigned((wire29 > ($signed(reg63) ^ "GThKM7k08slwZ"))));
            end
        end
      else
        begin
          if ("Ot8a5q39")
            begin
              reg46 = reg40;
              reg47 <= ({{(^(+reg56)),
                      wire32}} | $signed((-reg48[(1'h0):(1'h0)])));
              reg48 <= (8'h9f);
              reg50 = (reg61[(1'h0):(1'h0)] ?
                  (-$signed((reg63[(1'h0):(1'h0)] >>> (+(8'hb3))))) : $unsigned($signed((~|$signed(wire29)))));
            end
          else
            begin
              reg47 <= ($signed($unsigned(((~forvar46) <= ((8'haa) << reg47)))) ?
                  reg39[(3'h4):(3'h4)] : (-("tDL1O" ?
                      "" : {(forvar36 >> reg57)})));
              reg48 <= $signed(($unsigned($unsigned(reg63)) ?
                  $signed(forvar36[(1'h1):(1'h1)]) : (reg57 + (~&reg41[(4'ha):(3'h6)]))));
              reg50 = ($signed($unsigned((&(reg45 ?
                  reg47 : (8'hb7))))) ~^ $unsigned({$unsigned((reg43 ?
                      (8'hb8) : (8'h9d)))}));
              reg51 <= $unsigned((8'h9f));
            end
          for (forvar52 = (1'h0); (forvar52 < (3'h4)); forvar52 = (forvar52 + (1'h1)))
            begin
              reg53 <= reg55[(3'h4):(1'h1)];
              reg54 = $signed(($unsigned(((8'hb3) ? (+forvar46) : forvar54)) ?
                  $signed({(wire31 ? reg39 : reg38)}) : (wire30[(3'h4):(1'h0)] ?
                      reg40[(1'h0):(1'h0)] : (-wire30))));
            end
          reg55 <= wire32[(2'h3):(2'h3)];
          reg56 <= $signed((~$signed(reg60)));
          reg59 = ($unsigned($signed((!{wire29}))) | $unsigned({forvar36[(2'h3):(1'h1)],
              (~|(reg38 ? reg44 : reg58))}));
        end
    end
  module65 #() modinst168 (wire167, clk, wire31, reg57, reg55, reg45, wire28);
  assign wire169 = $unsigned(({($signed(reg47) | (reg53 != reg51)), reg39} ?
                       (8'ha4) : reg53[(3'h4):(2'h3)]));
  assign wire170 = (-((((reg55 == reg49) ?
                       (reg56 | reg56) : wire167[(1'h0):(1'h0)]) ^~ $unsigned($signed(reg52))) > (reg39[(3'h5):(2'h3)] ?
                       ($unsigned(wire31) ?
                           (reg58 ~^ reg35) : {wire31}) : reg57)));
  assign wire171 = ({wire31[(4'hf):(3'h7)]} <<< reg49);
  module172 #() modinst274 (wire273, clk, wire29, reg57, reg35, wire30);
  module275 #() modinst386 (wire385, clk, reg56, reg37, reg52, wire32, reg39);
  always
    @(posedge clk) begin
      if (reg55[(1'h0):(1'h0)])
        begin
          reg387 <= reg52[(3'h6):(3'h5)];
          reg388 = (reg63 > wire30);
          reg389 = (~((7'h42) >> (+((8'hac) ?
              $unsigned(reg37) : (^~wire169)))));
          for (forvar390 = (1'h0); (forvar390 < (2'h3)); forvar390 = (forvar390 + (1'h1)))
            begin
              reg391 = $signed(wire30);
              reg392 = wire171;
              reg393 <= ({$unsigned(((reg51 && wire169) & (reg35 | reg35))),
                  ($signed((&wire385)) | reg57[(4'h9):(4'h8)])} && $signed(wire169));
              reg394 = reg393[(3'h6):(1'h0)];
              reg395 <= reg52[(2'h3):(2'h3)];
            end
          reg396 = $unsigned((!($signed((reg45 << reg51)) << wire169[(3'h5):(3'h4)])));
        end
      else
        begin
          for (forvar387 = (1'h0); (forvar387 < (1'h0)); forvar387 = (forvar387 + (1'h1)))
            begin
              reg390 <= "SuJ2fsv32TWAoM0Toxn";
              reg391 = (reg390 ?
                  {$signed(reg396), "pA5"} : ($unsigned(({(8'hb8)} ?
                      (reg396 ? (8'hb6) : (8'hbc)) : ((8'hbe) ?
                          reg389 : forvar387))) <= (~|(((8'hb2) >= reg62) ?
                      ((8'ha5) && reg39) : wire171[(3'h7):(3'h6)]))));
            end
          for (forvar392 = (1'h0); (forvar392 < (1'h1)); forvar392 = (forvar392 + (1'h1)))
            begin
              reg394 = $signed({$unsigned(($unsigned(reg52) >>> (reg48 > reg387)))});
              reg395 <= (!(8'hb7));
              reg396 = ((~|reg56) & "72qdMAJpv2ZMDbvDpGh");
            end
          for (forvar397 = (1'h0); (forvar397 < (2'h2)); forvar397 = (forvar397 + (1'h1)))
            begin
              reg398 = (^~reg57[(1'h0):(1'h0)]);
              reg399 <= forvar397;
            end
          reg400 <= (^~reg47);
          reg401 <= $unsigned((({$signed(reg394)} != $unsigned($signed(reg56))) ?
              {reg396} : ((&wire385) ?
                  (reg394[(3'h4):(3'h4)] == (!reg392)) : (~(-reg393)))));
        end
      reg402 <= $signed((((((8'ha0) != wire30) <<< reg35) ?
          reg393[(3'h4):(1'h1)] : {wire169}) ^ reg398[(3'h5):(1'h1)]));
      for (forvar403 = (1'h0); (forvar403 < (3'h4)); forvar403 = (forvar403 + (1'h1)))
        begin
          for (forvar404 = (1'h0); (forvar404 < (3'h4)); forvar404 = (forvar404 + (1'h1)))
            begin
              reg405 <= {(reg400[(1'h1):(1'h0)] ? {(-reg393)} : reg391),
                  $signed((reg396[(1'h1):(1'h1)] < $signed((wire169 ?
                      (8'ha4) : reg48))))};
              reg406 = ($signed($signed({(reg45 <= reg390),
                      {wire32, wire30}})) ?
                  (^~reg57) : $unsigned({($signed(wire30) + (reg47 ?
                          reg387 : wire28)),
                      (reg390[(4'ha):(3'h5)] ?
                          $signed(reg45) : (reg39 ~^ reg391))}));
            end
        end
    end
  assign wire407 = wire28[(4'hd):(2'h2)];
  assign wire408 = (8'hbc);
  module409 #() modinst472 (.wire414(wire169), .wire413(wire385), .wire411(reg402), .clk(clk), .wire410(reg48), .y(wire471), .wire412(reg51));
  assign wire473 = wire385;
  assign wire474 = (wire171 >> ({(reg53[(3'h6):(3'h6)] ?
                           reg45[(1'h0):(1'h0)] : $unsigned(reg57)),
                       wire31} > (reg58 ?
                       ("Rcf8lD1EVAvc3KpRLOs" * (-wire385)) : ($unsigned((8'ha6)) ?
                           reg400[(4'hb):(3'h7)] : (^~reg63)))));
  assign wire475 = reg401[(4'he):(2'h2)];
  assign wire476 = {(reg387 + (&{(8'hb4)}))};
  module477 #() modinst584 (wire583, clk, reg405, wire273, reg58, reg401);
  always
    @(posedge clk) begin
      for (forvar585 = (1'h0); (forvar585 < (2'h2)); forvar585 = (forvar585 + (1'h1)))
        begin
          for (forvar586 = (1'h0); (forvar586 < (3'h4)); forvar586 = (forvar586 + (1'h1)))
            begin
              reg587 = ((reg37 ?
                  reg55[(4'hf):(4'h9)] : reg39[(1'h1):(1'h1)]) >>> ((~wire471) - $signed(($unsigned(wire171) ?
                  (reg390 >>> reg387) : "IXGPHQrSwR4om"))));
            end
        end
      for (forvar588 = (1'h0); (forvar588 < (1'h0)); forvar588 = (forvar588 + (1'h1)))
        begin
          if ($signed($signed((reg399[(5'h10):(3'h6)] != $signed((reg387 ?
              reg390 : wire407))))))
            begin
              reg589 = reg387;
              reg590 = (reg45 ? (7'h44) : wire31[(3'h6):(1'h0)]);
              reg591 <= {$unsigned({{(|reg49), (8'hbd)}}),
                  ($signed(reg590) - $unsigned(($unsigned(reg390) ?
                      "QAnM" : $signed(reg399))))};
              reg592 <= {$signed(reg399[(4'hc):(4'hc)])};
              reg593 <= ($unsigned(reg45[(3'h5):(3'h4)]) ?
                  wire169[(4'h8):(2'h2)] : ((~|$signed((&wire170))) ?
                      reg399 : (!(reg63[(2'h2):(1'h1)] | (reg39 ?
                          reg591 : wire28)))));
            end
          else
            begin
              reg589 = $signed((8'hab));
              reg591 <= $signed($signed($unsigned($unsigned(reg589))));
              reg594 = $signed(((reg48[(2'h3):(2'h3)] ?
                      wire29 : $signed(((8'ha4) ? reg53 : reg400))) ?
                  ((&(reg592 ? wire473 : (8'ha9))) & (wire29 ?
                      $signed((8'hbd)) : {reg405,
                          reg395})) : $unsigned($unsigned(((8'ha6) & forvar586)))));
              reg595 <= "AoSLhNuEs3emQMDI9";
              reg596 <= (reg395[(4'ha):(1'h1)] ?
                  ((($unsigned((8'ha7)) ?
                      wire407 : $unsigned((7'h41))) >> (reg45[(1'h0):(1'h0)] ?
                      (reg402 != (8'ha0)) : $signed(wire471))) == $unsigned($unsigned((reg55 == forvar588)))) : $signed($unsigned(("nZpssOo" ^ wire167[(4'h8):(1'h0)]))));
            end
          for (forvar597 = (1'h0); (forvar597 < (1'h1)); forvar597 = (forvar597 + (1'h1)))
            begin
              reg598 = "1No85ee1us";
              reg599 = (7'h42);
              reg600 <= $signed((|(((~^(8'ha2)) ? wire28 : $unsigned(wire171)) ?
                  wire476[(1'h1):(1'h1)] : ($unsigned(reg595) & (reg593 ?
                      (8'ha6) : reg37)))));
              reg601 = $unsigned(forvar585[(4'he):(4'hc)]);
              reg602 <= (~&$signed($signed(wire29)));
            end
          reg603 = $unsigned("NWmNScFRwoYUXLoOD4XQ");
        end
      reg604 <= reg39;
      if ((8'hbc))
        begin
          reg605 <= (8'ha1);
          for (forvar606 = (1'h0); (forvar606 < (2'h3)); forvar606 = (forvar606 + (1'h1)))
            begin
              reg607 <= $signed(forvar606);
              reg608 <= ({({wire474[(2'h2):(1'h1)]} > ($unsigned(wire32) ^~ (wire407 ?
                      (8'hb7) : reg590)))} - $signed(($unsigned($unsigned(reg53)) ?
                  $signed({wire476, (8'hb7)}) : $signed($unsigned(reg52)))));
            end
        end
      else
        begin
          reg606 = ($unsigned(reg608[(4'he):(1'h0)]) << $signed((reg589 ?
              ((reg401 ^ wire475) ?
                  ((8'ha4) * reg45) : $unsigned(reg592)) : (~^reg402[(4'h8):(4'h8)]))));
          reg607 <= (wire473[(4'h8):(1'h0)] * wire171);
          reg608 <= $signed(wire170);
          if (reg387)
            begin
              reg609 = $signed((reg402[(5'h14):(5'h11)] < ($unsigned(reg605[(3'h5):(3'h4)]) ?
                  (-(|reg599)) : {(forvar606 ? reg51 : wire171), (~&reg600)})));
              reg610 = ($unsigned((7'h43)) & "R2iCao");
              reg611 = $signed($unsigned($unsigned(reg405)));
              reg612 <= wire407;
              reg613 <= (reg593[(1'h1):(1'h1)] ?
                  $unsigned((|((reg62 ? reg57 : wire407) ?
                      {reg590} : {(8'hac)}))) : $unsigned(reg610));
            end
          else
            begin
              reg609 = (wire476 * $unsigned($unsigned($signed(reg593))));
              reg612 <= (~^reg35);
            end
          for (forvar614 = (1'h0); (forvar614 < (1'h1)); forvar614 = (forvar614 + (1'h1)))
            begin
              reg615 = forvar614[(3'h7):(2'h2)];
              reg616 <= reg599[(2'h2):(2'h2)];
              reg617 <= (+$signed(reg611[(4'ha):(4'ha)]));
            end
        end
      for (forvar618 = (1'h0); (forvar618 < (1'h1)); forvar618 = (forvar618 + (1'h1)))
        begin
          for (forvar619 = (1'h0); (forvar619 < (3'h4)); forvar619 = (forvar619 + (1'h1)))
            begin
              reg620 = (~|(^~reg608[(4'hc):(4'ha)]));
              reg621 = (reg595[(4'h8):(2'h3)] ?
                  $unsigned($signed((^$unsigned(reg387)))) : (~&(~&((~|reg400) + $unsigned((8'h9c))))));
              reg622 = $unsigned(({($unsigned(reg35) < reg53[(3'h7):(2'h2)]),
                  ($signed(reg47) ?
                      (reg609 ?
                          wire583 : wire28) : (7'h41))} < (wire28[(1'h1):(1'h1)] >= ((reg607 != reg615) ?
                  $signed(reg49) : reg587))));
              reg623 = forvar618[(4'h8):(3'h5)];
            end
          if ($unsigned(($unsigned($unsigned($unsigned(wire170))) ^~ (((^~reg400) ?
              (~forvar597) : $signed(wire385)) & reg587))))
            begin
              reg624 = reg595;
              reg625 <= (-wire273);
              reg626 <= wire30[(3'h4):(2'h3)];
              reg627 <= {{(($unsigned(wire32) >> (!wire471)) >= $signed($signed(reg623))),
                      ($signed(wire385) ? reg56[(4'he):(4'hb)] : reg48)}};
              reg628 = "";
            end
          else
            begin
              reg625 <= $signed((!reg390[(1'h1):(1'h0)]));
              reg628 = $signed($signed($signed(((reg53 ? reg395 : reg387) ?
                  reg53[(5'h10):(4'h8)] : wire29))));
            end
          if ((^$signed((reg613[(2'h3):(2'h2)] ? $signed(wire170) : reg612))))
            begin
              reg629 <= $unsigned((~$unsigned($unsigned((!wire171)))));
              reg630 = $unsigned(wire474);
              reg631 = (reg405[(3'h5):(2'h3)] ?
                  $unsigned($unsigned(((reg605 ?
                      (8'h9e) : reg612) * forvar618))) : {wire170,
                      reg402[(5'h15):(3'h4)]});
              reg632 = $unsigned($unsigned(wire475));
              reg633 = (8'hbf);
            end
          else
            begin
              reg629 <= (^~(~|{(&(reg608 ? forvar618 : reg632))}));
              reg634 <= $unsigned({(~|wire170)});
              reg635 <= ((wire385 ?
                      ($unsigned(((8'hb4) ? reg399 : wire475)) ?
                          $signed((8'hb6)) : forvar585) : wire28[(5'h10):(4'hb)]) ?
                  (reg611 == $signed(reg62)) : ((($unsigned(forvar618) ?
                      reg48[(4'h8):(3'h7)] : ((8'haa) <<< (8'hbd))) - reg37[(4'h8):(1'h1)]) >> ($signed({reg590}) || $signed((wire583 << wire169)))));
              reg636 <= reg623[(4'hc):(1'h0)];
            end
          reg637 <= ($unsigned((reg623[(5'h10):(1'h0)] | $signed((wire28 ?
              reg387 : forvar618)))) * $signed(($unsigned(((8'ha3) != (8'hbe))) <<< (reg628 ?
              (reg594 ? reg47 : reg51) : forvar619))));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module477
#(parameter param581 = ((~|(|(((7'h42) ? (7'h40) : (7'h42)) ^ ((8'h9c) ? (7'h41) : (8'ha9))))) ? ({(|{(8'hba)}), {((8'hae) || (8'ha2)), (8'hbd)}} ? ((((8'h9d) >>> (8'ha0)) <= ((8'hb8) == (8'hb3))) ? (((7'h44) >> (8'h9e)) ~^ ((8'ha4) ? (8'ha4) : (8'ha9))) : ((^(8'ha0)) ? (~|(7'h43)) : {(8'ha2)})) : (((8'hab) & ((8'hb2) & (8'ha7))) ? ((~^(8'haa)) ? ((8'h9d) ? (8'hb3) : (8'hb7)) : ((8'ha7) <= (8'ha7))) : (^{(8'h9e), (8'ha5)}))) : ((~({(8'hbe), (8'hb8)} || (8'hb5))) ^~ (({(8'hb1), (8'hac)} ? ((8'h9e) * (8'ha0)) : ((8'ha0) != (8'hb7))) >>> (-(~|(8'haa)))))), 
parameter param582 = ((-(~|(|param581))) <= (^~{(8'hbc)})))
(y, clk, wire481, wire480, wire479, wire478);
  output wire [(32'h48e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire481;
  input wire [(5'h11):(1'h0)] wire480;
  input wire signed [(4'h8):(1'h0)] wire479;
  input wire signed [(2'h3):(1'h0)] wire478;
  wire [(3'h7):(1'h0)] wire580;
  wire [(4'h9):(1'h0)] wire579;
  wire [(2'h3):(1'h0)] wire578;
  wire signed [(5'h14):(1'h0)] wire577;
  wire signed [(4'hc):(1'h0)] wire576;
  reg [(4'hd):(1'h0)] reg575 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg574 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg570 = (1'h0);
  reg [(4'h8):(1'h0)] reg569 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg568 = (1'h0);
  reg [(4'ha):(1'h0)] reg567 = (1'h0);
  reg [(4'he):(1'h0)] reg566 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg565 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg563 = (1'h0);
  reg [(2'h3):(1'h0)] reg561 = (1'h0);
  reg [(4'hc):(1'h0)] reg559 = (1'h0);
  reg [(4'ha):(1'h0)] reg557 = (1'h0);
  reg [(3'h7):(1'h0)] reg555 = (1'h0);
  reg [(5'h15):(1'h0)] reg551 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg552 = (1'h0);
  reg [(5'h15):(1'h0)] reg550 = (1'h0);
  reg [(5'h12):(1'h0)] reg549 = (1'h0);
  reg [(2'h2):(1'h0)] reg548 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg545 = (1'h0);
  reg [(5'h15):(1'h0)] reg542 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg541 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg540 = (1'h0);
  reg [(4'he):(1'h0)] reg537 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg530 = (1'h0);
  reg [(4'hf):(1'h0)] reg529 = (1'h0);
  reg [(2'h3):(1'h0)] reg528 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg526 = (1'h0);
  reg [(5'h10):(1'h0)] reg525 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg524 = (1'h0);
  reg [(3'h7):(1'h0)] reg523 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg514 = (1'h0);
  reg [(4'h9):(1'h0)] reg510 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg520 = (1'h0);
  reg [(4'hd):(1'h0)] reg519 = (1'h0);
  reg [(3'h7):(1'h0)] reg516 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg513 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg509 = (1'h0);
  reg [(5'h14):(1'h0)] reg508 = (1'h0);
  reg [(5'h11):(1'h0)] reg504 = (1'h0);
  reg [(4'ha):(1'h0)] reg503 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg502 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg501 = (1'h0);
  reg [(5'h14):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg498 = (1'h0);
  reg [(2'h3):(1'h0)] reg497 = (1'h0);
  reg [(5'h15):(1'h0)] reg493 = (1'h0);
  reg [(2'h2):(1'h0)] reg492 = (1'h0);
  reg [(4'hc):(1'h0)] reg489 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg485 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg483 = (1'h0);
  reg [(4'ha):(1'h0)] reg573 = (1'h0);
  reg [(4'hf):(1'h0)] reg572 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg571 = (1'h0);
  reg [(3'h4):(1'h0)] forvar564 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg562 = (1'h0);
  reg [(2'h3):(1'h0)] reg560 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar558 = (1'h0);
  reg [(4'hd):(1'h0)] reg556 = (1'h0);
  reg [(4'hd):(1'h0)] reg554 = (1'h0);
  reg signed [(4'he):(1'h0)] reg553 = (1'h0);
  reg [(5'h10):(1'h0)] forvar551 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg547 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar546 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg544 = (1'h0);
  reg [(4'hf):(1'h0)] reg543 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg539 = (1'h0);
  reg [(3'h6):(1'h0)] forvar538 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg536 = (1'h0);
  reg [(4'he):(1'h0)] reg535 = (1'h0);
  reg [(4'he):(1'h0)] reg534 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar533 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg532 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg531 = (1'h0);
  reg [(4'hb):(1'h0)] forvar527 = (1'h0);
  reg [(2'h3):(1'h0)] reg527 = (1'h0);
  reg [(3'h6):(1'h0)] reg522 = (1'h0);
  reg [(4'h9):(1'h0)] forvar511 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg521 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg518 = (1'h0);
  reg [(4'he):(1'h0)] reg517 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg515 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar514 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg512 = (1'h0);
  reg [(4'hf):(1'h0)] reg511 = (1'h0);
  reg [(5'h14):(1'h0)] forvar510 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg507 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar506 = (1'h0);
  reg [(3'h4):(1'h0)] reg505 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg500 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg496 = (1'h0);
  reg [(5'h14):(1'h0)] forvar495 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg494 = (1'h0);
  reg [(3'h5):(1'h0)] reg491 = (1'h0);
  reg [(4'h8):(1'h0)] forvar490 = (1'h0);
  reg [(4'h9):(1'h0)] reg488 = (1'h0);
  reg [(4'h8):(1'h0)] forvar487 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg486 = (1'h0);
  reg [(4'hc):(1'h0)] forvar484 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar482 = (1'h0);
  assign y = {wire580,
                 wire579,
                 wire578,
                 wire577,
                 wire576,
                 reg575,
                 reg574,
                 reg570,
                 reg569,
                 reg568,
                 reg567,
                 reg566,
                 reg565,
                 reg563,
                 reg561,
                 reg559,
                 reg557,
                 reg555,
                 reg551,
                 reg552,
                 reg550,
                 reg549,
                 reg548,
                 reg545,
                 reg542,
                 reg541,
                 reg540,
                 reg537,
                 reg530,
                 reg529,
                 reg528,
                 reg526,
                 reg525,
                 reg524,
                 reg523,
                 reg514,
                 reg510,
                 reg520,
                 reg519,
                 reg516,
                 reg513,
                 reg509,
                 reg508,
                 reg504,
                 reg503,
                 reg502,
                 reg501,
                 reg499,
                 reg498,
                 reg497,
                 reg493,
                 reg492,
                 reg489,
                 reg485,
                 reg483,
                 reg573,
                 reg572,
                 reg571,
                 forvar564,
                 reg562,
                 reg560,
                 forvar558,
                 reg556,
                 reg554,
                 reg553,
                 forvar551,
                 reg547,
                 forvar546,
                 reg544,
                 reg543,
                 reg539,
                 forvar538,
                 reg536,
                 reg535,
                 reg534,
                 forvar533,
                 reg532,
                 reg531,
                 forvar527,
                 reg527,
                 reg522,
                 forvar511,
                 reg521,
                 reg518,
                 reg517,
                 reg515,
                 forvar514,
                 reg512,
                 reg511,
                 forvar510,
                 reg507,
                 forvar506,
                 reg505,
                 reg500,
                 reg496,
                 forvar495,
                 reg494,
                 reg491,
                 forvar490,
                 reg488,
                 forvar487,
                 reg486,
                 forvar484,
                 forvar482,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar482 = (1'h0); (forvar482 < (3'h4)); forvar482 = (forvar482 + (1'h1)))
        begin
          reg483 <= wire480[(2'h3):(2'h3)];
          for (forvar484 = (1'h0); (forvar484 < (3'h4)); forvar484 = (forvar484 + (1'h1)))
            begin
              reg485 <= {{$unsigned($unsigned(reg483)),
                      $unsigned(((~|forvar482) ?
                          $signed(forvar482) : (reg483 >>> wire481)))}};
              reg486 = $signed($unsigned(wire478));
            end
          for (forvar487 = (1'h0); (forvar487 < (2'h3)); forvar487 = (forvar487 + (1'h1)))
            begin
              reg488 = (forvar484 ?
                  $unsigned($unsigned($signed((forvar482 * wire479)))) : forvar487[(1'h1):(1'h0)]);
              reg489 <= (~(reg483 ~^ wire478[(1'h1):(1'h0)]));
            end
          for (forvar490 = (1'h0); (forvar490 < (1'h1)); forvar490 = (forvar490 + (1'h1)))
            begin
              reg491 = ((forvar487[(1'h0):(1'h0)] ?
                      ("bUTSWHn2MH" ?
                          reg489[(3'h4):(1'h1)] : (forvar490 - (~wire478))) : (("8WrvHtsfz5NqLRy" < forvar484) ?
                          $signed((!forvar484)) : (^~(forvar487 != forvar482)))) ?
                  $signed($unsigned(((forvar482 ?
                      forvar490 : wire480) - (&(8'hb0))))) : {(($unsigned(reg486) ?
                          $signed(reg485) : $unsigned(forvar490)) >>> (8'hab)),
                      {$unsigned({(8'hbc)}), forvar490[(3'h5):(2'h3)]}});
              reg492 <= reg483[(4'h9):(1'h0)];
              reg493 <= {(8'ha6), (-$unsigned(wire479[(1'h0):(1'h0)]))};
              reg494 = wire480;
            end
        end
      for (forvar495 = (1'h0); (forvar495 < (2'h3)); forvar495 = (forvar495 + (1'h1)))
        begin
          reg496 = ((8'ha5) * $unsigned((wire480 | ((reg494 >= reg485) << reg494))));
          reg497 <= $signed((~^({"gGhH"} ?
              (^~(reg485 ? reg483 : forvar490)) : {reg485,
                  ((8'ha8) | (7'h41))})));
          if ($signed((8'hb6)))
            begin
              reg498 <= ($signed((8'hbd)) & (!{{((8'ha4) * wire481)},
                  (~|$signed(wire481))}));
              reg499 <= reg489;
              reg500 = reg496;
              reg501 <= (7'h43);
            end
          else
            begin
              reg498 <= reg483[(5'h12):(4'hf)];
              reg500 = $unsigned($unsigned(reg488[(3'h6):(1'h0)]));
              reg501 <= reg497;
              reg502 <= $unsigned(($unsigned($signed($signed(forvar495))) <= reg499[(4'he):(4'hb)]));
              reg503 <= $unsigned($unsigned(wire478));
            end
        end
      if ($unsigned((8'hb5)))
        begin
          reg504 <= {$unsigned(reg483[(3'h4):(1'h1)])};
        end
      else
        begin
          reg505 = $signed((^reg501[(4'hf):(4'hc)]));
          for (forvar506 = (1'h0); (forvar506 < (3'h4)); forvar506 = (forvar506 + (1'h1)))
            begin
              reg507 = ({(((~|reg493) + {reg486}) ?
                          reg489[(1'h1):(1'h0)] : $signed((reg492 ?
                              (8'hb9) : (8'h9f))))} ?
                  reg504[(2'h2):(1'h1)] : reg492[(1'h1):(1'h0)]);
              reg508 <= (($signed(wire479) ?
                  ((~|(reg502 || forvar482)) * (|(+reg489))) : (((7'h41) ?
                      ((8'hbb) & reg504) : (forvar495 >> reg496)) ^ (^~reg488[(3'h7):(3'h4)]))) | (8'h9c));
              reg509 <= (^($unsigned({(~|(7'h40))}) ?
                  (~^((reg500 ?
                      (8'ha0) : forvar495) || (8'hb0))) : ($unsigned((wire481 ?
                      reg503 : reg492)) < ((reg502 - forvar490) ?
                      (reg486 != reg503) : (wire480 ? reg501 : wire478)))));
            end
        end
      if ($unsigned($unsigned({{reg504}, (|(forvar490 ? reg509 : reg504))})))
        begin
          for (forvar510 = (1'h0); (forvar510 < (2'h3)); forvar510 = (forvar510 + (1'h1)))
            begin
              reg511 = ({wire479[(1'h0):(1'h0)],
                      $signed($unsigned({forvar484}))} ?
                  {(reg489[(4'h9):(4'h9)] >>> {(reg485 ? wire480 : forvar482),
                          (forvar506 ? reg504 : reg499)}),
                      ($unsigned((reg493 ? reg483 : reg498)) ?
                          (!$unsigned(reg488)) : (~^reg497))} : $unsigned((((^reg488) ?
                      reg501[(4'h9):(2'h3)] : forvar495[(5'h13):(1'h1)]) == $signed({forvar484}))));
              reg512 = reg483[(4'he):(1'h0)];
              reg513 <= (-$signed((reg504[(4'hf):(1'h0)] ?
                  (&(reg494 == reg498)) : $signed(((8'hb5) == forvar484)))));
            end
          for (forvar514 = (1'h0); (forvar514 < (1'h1)); forvar514 = (forvar514 + (1'h1)))
            begin
              reg515 = $unsigned(reg497[(2'h3):(1'h0)]);
              reg516 <= $unsigned((+(~&((&forvar484) ?
                  (reg504 ? reg512 : (8'haf)) : (forvar506 ?
                      reg507 : (8'hb6))))));
              reg517 = forvar495;
            end
          if ({reg486[(4'ha):(3'h6)], $unsigned({reg497[(2'h2):(1'h0)]})})
            begin
              reg518 = forvar506;
              reg519 <= $unsigned($unsigned((|(8'hb7))));
              reg520 <= wire479[(4'h8):(1'h1)];
            end
          else
            begin
              reg519 <= reg505;
              reg521 = $unsigned({(reg498 ?
                      ((&reg496) ?
                          reg497 : $unsigned((8'ha6))) : forvar490[(3'h4):(1'h1)]),
                  (+{(reg507 || reg488), (reg509 ^ forvar514)})});
            end
        end
      else
        begin
          reg510 <= "ckqiOcO";
          for (forvar511 = (1'h0); (forvar511 < (1'h1)); forvar511 = (forvar511 + (1'h1)))
            begin
              reg512 = reg517;
              reg513 <= reg512[(3'h4):(2'h3)];
              reg514 <= reg497;
              reg516 <= ($unsigned($unsigned(wire479)) ?
                  (!((((8'hb6) ? reg503 : reg509) ?
                          (reg505 ^~ forvar490) : $unsigned(forvar490)) ?
                      forvar514 : reg496[(3'h4):(2'h3)])) : reg499[(5'h12):(4'h9)]);
              reg519 <= (+"oFBwuVXD");
            end
          if ({$unsigned((~forvar506[(3'h7):(3'h7)])),
              $unsigned(($unsigned((reg488 ?
                  forvar487 : reg512)) >>> forvar511[(4'h9):(2'h3)]))})
            begin
              reg521 = $signed("yb0msILVpz");
              reg522 = $signed($unsigned(reg488));
              reg523 <= reg483[(3'h6):(1'h1)];
              reg524 <= reg497;
            end
          else
            begin
              reg520 <= ($signed(reg507[(3'h4):(2'h2)]) > forvar510[(4'h9):(3'h5)]);
              reg521 = forvar514;
              reg523 <= reg514;
            end
          reg525 <= {(~^(~^$unsigned(reg511[(4'he):(4'hc)])))};
          reg526 <= (^~reg505[(3'h4):(3'h4)]);
        end
      if (reg489)
        begin
          reg527 = reg505[(1'h1):(1'h1)];
        end
      else
        begin
          for (forvar527 = (1'h0); (forvar527 < (1'h0)); forvar527 = (forvar527 + (1'h1)))
            begin
              reg528 <= $signed(forvar506);
              reg529 <= reg521[(2'h2):(1'h0)];
              reg530 <= $unsigned((^~("g3ziFVE" & reg500)));
              reg531 = $unsigned(wire479[(2'h3):(2'h3)]);
            end
          reg532 = $signed("12utbuvbvCHm3y5");
          for (forvar533 = (1'h0); (forvar533 < (1'h0)); forvar533 = (forvar533 + (1'h1)))
            begin
              reg534 = ($unsigned(reg499[(4'hd):(1'h1)]) ?
                  reg491[(2'h2):(1'h0)] : (7'h43));
              reg535 = ((reg498[(3'h4):(1'h0)] || forvar514) ? reg485 : reg534);
              reg536 = $signed(reg524[(4'h9):(1'h0)]);
              reg537 <= forvar527[(3'h7):(3'h6)];
            end
          for (forvar538 = (1'h0); (forvar538 < (2'h2)); forvar538 = (forvar538 + (1'h1)))
            begin
              reg539 = reg507;
            end
          reg540 <= ((~^$unsigned($unsigned(reg516[(3'h4):(2'h3)]))) ?
              reg530[(1'h1):(1'h1)] : $signed($unsigned($unsigned((reg536 ?
                  reg492 : reg522)))));
        end
    end
  always
    @(posedge clk) begin
      if ($signed($signed(reg499)))
        begin
          reg541 <= reg514;
          reg542 <= reg520;
          reg543 = $unsigned(({{reg529[(2'h3):(2'h2)], (~|reg523)},
                  wire479[(2'h2):(1'h0)]} ?
              ((reg513 || (!wire478)) << ((8'ha4) | (7'h43))) : "FzC"));
        end
      else
        begin
          reg541 <= wire478;
          if ({reg493,
              ((((reg493 ? reg520 : (8'hba)) ?
                      reg492[(2'h2):(2'h2)] : ((8'ha2) <<< wire478)) > $signed({reg510})) ?
                  wire481 : $signed((reg492[(1'h0):(1'h0)] && (reg525 ~^ reg520))))})
            begin
              reg543 = (8'hab);
            end
          else
            begin
              reg542 <= $signed(reg508);
              reg543 = (~^$unsigned({wire480[(3'h7):(3'h7)]}));
              reg544 = {$signed({reg526, (8'hb6)})};
              reg545 <= $signed(reg483[(4'he):(3'h4)]);
            end
          for (forvar546 = (1'h0); (forvar546 < (1'h1)); forvar546 = (forvar546 + (1'h1)))
            begin
              reg547 = (($unsigned($signed($unsigned(reg544))) & (reg510 ?
                  (+$unsigned(reg526)) : ($signed(reg542) == $signed(reg502)))) && "0JNuhR8LCQ");
              reg548 <= ((~|{"EDVdyr3u0lv44aXL"}) < ((~|{wire481,
                  (8'hbb)}) | (8'hb4)));
              reg549 <= $signed(($signed($unsigned($signed(reg502))) ?
                  ((+(8'h9f)) ~^ $signed((8'hbf))) : ((wire479 <= (reg514 >> reg519)) ?
                      (8'hbd) : reg498[(1'h0):(1'h0)])));
            end
          reg550 <= ({$signed(reg508[(4'h8):(3'h7)])} ?
              ($unsigned(reg545) ?
                  $signed((reg547[(2'h2):(1'h1)] ~^ reg483[(4'hb):(2'h3)])) : ($signed((reg549 >> reg526)) ?
                      (reg497 ?
                          {reg525} : (reg502 || wire478)) : ({reg525} + $unsigned(reg525)))) : $signed($signed($signed("l"))));
        end
      if ((-{$unsigned(($unsigned(reg524) ?
              ((7'h41) ? reg501 : (7'h43)) : reg537))}))
        begin
          for (forvar551 = (1'h0); (forvar551 < (3'h4)); forvar551 = (forvar551 + (1'h1)))
            begin
              reg552 <= reg503[(3'h4):(2'h3)];
            end
        end
      else
        begin
          if ($signed((~^reg552)))
            begin
              reg551 <= (+"pNRLFeTbnDE5I2MwxA0");
            end
          else
            begin
              reg553 = $unsigned(reg497);
              reg554 = wire479[(1'h0):(1'h0)];
              reg555 <= ((~(~$signed((~reg553)))) <= ((-(+reg525[(4'he):(3'h7)])) ~^ (reg544[(4'hd):(2'h2)] || (!reg544[(3'h4):(1'h0)]))));
              reg556 = (^reg508);
            end
          reg557 <= (-(reg503[(1'h1):(1'h0)] <= ($signed((^~reg548)) ?
              reg510 : (8'hbf))));
        end
      if ($signed($unsigned((~&{{reg550}, (reg516 ? reg523 : reg524)}))))
        begin
          for (forvar558 = (1'h0); (forvar558 < (1'h0)); forvar558 = (forvar558 + (1'h1)))
            begin
              reg559 <= (reg550 ^ reg502);
              reg560 = reg523[(1'h1):(1'h1)];
              reg561 <= $signed($signed(reg528[(1'h1):(1'h1)]));
              reg562 = reg489;
            end
        end
      else
        begin
          for (forvar558 = (1'h0); (forvar558 < (2'h3)); forvar558 = (forvar558 + (1'h1)))
            begin
              reg560 = (($signed((((8'hbf) ? reg502 : reg540) ?
                      $unsigned(reg483) : (8'hb4))) ?
                  (|$unsigned(wire478[(2'h2):(2'h2)])) : $signed((reg523 || (reg559 ?
                      (7'h40) : forvar558)))) != {{(-(reg483 ?
                          reg483 : (8'hae))),
                      reg516},
                  reg552[(2'h3):(2'h2)]});
              reg561 <= reg549[(4'h8):(3'h6)];
              reg563 <= reg550[(4'h8):(1'h1)];
            end
          for (forvar564 = (1'h0); (forvar564 < (1'h0)); forvar564 = (forvar564 + (1'h1)))
            begin
              reg565 <= reg503;
              reg566 <= {$unsigned(reg562[(4'h9):(3'h6)]),
                  $unsigned({$signed("VzoLQ30LyhZpEXx"), (^(!(8'hb7)))})};
              reg567 <= reg509;
              reg568 <= reg513;
              reg569 <= {reg497[(2'h3):(1'h0)]};
            end
          reg570 <= $unsigned((^~(("vxLJhxBB7" ?
              (8'hb1) : {reg540, reg551}) != "9EMUZASsKk")));
          reg571 = (~forvar546);
          if ($unsigned((reg553[(3'h6):(2'h2)] > $unsigned($unsigned((reg544 ?
              reg559 : reg513))))))
            begin
              reg572 = {reg560,
                  (("ylDsBf" | ((reg545 * reg485) >> reg542[(5'h11):(4'h8)])) ?
                      $signed($unsigned("KxAnPFiX5xXILJLM")) : {$signed((reg524 ~^ reg510)),
                          $unsigned((-reg499))})};
            end
          else
            begin
              reg572 = reg497;
              reg573 = reg568;
              reg574 <= reg548;
            end
        end
      reg575 <= ($unsigned(reg568[(3'h5):(1'h1)]) < {reg555});
    end
  assign wire576 = $signed((reg503[(3'h5):(2'h2)] ? {reg514, reg519} : reg499));
  assign wire577 = (^reg537);
  assign wire578 = ($unsigned((^~{(!reg526), reg525[(4'h8):(3'h4)]})) ?
                       ($unsigned((|((8'haa) ?
                           (8'h9d) : wire481))) <<< $signed($unsigned($unsigned(reg570)))) : reg548[(2'h2):(2'h2)]);
  assign wire579 = reg489[(4'hb):(4'h8)];
  assign wire580 = $unsigned(($unsigned(reg565[(2'h3):(1'h0)]) ?
                       ({$signed(wire481)} ?
                           (~^reg541) : $unsigned((^~wire481))) : (reg557 || $signed((reg540 >= (8'ha9))))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module409
#(parameter param470 = (7'h40))
(y, clk, wire414, wire413, wire412, wire411, wire410);
  output wire [(32'h2b3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire414;
  input wire signed [(5'h14):(1'h0)] wire413;
  input wire [(5'h12):(1'h0)] wire412;
  input wire [(4'hb):(1'h0)] wire411;
  input wire [(4'h9):(1'h0)] wire410;
  wire [(4'h8):(1'h0)] wire469;
  wire [(4'hd):(1'h0)] wire468;
  wire signed [(5'h13):(1'h0)] wire416;
  wire signed [(4'ha):(1'h0)] wire415;
  reg signed [(4'hc):(1'h0)] reg467 = (1'h0);
  reg signed [(4'he):(1'h0)] reg465 = (1'h0);
  reg [(5'h11):(1'h0)] reg463 = (1'h0);
  reg [(4'h8):(1'h0)] reg462 = (1'h0);
  reg [(5'h13):(1'h0)] reg458 = (1'h0);
  reg [(5'h13):(1'h0)] reg457 = (1'h0);
  reg [(5'h15):(1'h0)] reg455 = (1'h0);
  reg [(5'h15):(1'h0)] reg454 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg452 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg451 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg450 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg444 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg442 = (1'h0);
  reg [(4'he):(1'h0)] reg441 = (1'h0);
  reg [(5'h11):(1'h0)] reg436 = (1'h0);
  reg [(4'ha):(1'h0)] reg433 = (1'h0);
  reg [(5'h10):(1'h0)] reg432 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg430 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg421 = (1'h0);
  reg [(3'h6):(1'h0)] reg426 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg425 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg424 = (1'h0);
  reg [(3'h6):(1'h0)] reg423 = (1'h0);
  reg signed [(4'he):(1'h0)] reg422 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg419 = (1'h0);
  reg [(4'hc):(1'h0)] reg418 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg466 = (1'h0);
  reg [(3'h7):(1'h0)] reg464 = (1'h0);
  reg [(5'h12):(1'h0)] reg461 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg460 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg459 = (1'h0);
  reg [(3'h6):(1'h0)] reg456 = (1'h0);
  reg [(4'hc):(1'h0)] reg453 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar449 = (1'h0);
  reg [(3'h7):(1'h0)] reg448 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg447 = (1'h0);
  reg [(5'h10):(1'h0)] reg446 = (1'h0);
  reg [(4'hc):(1'h0)] reg445 = (1'h0);
  reg [(3'h4):(1'h0)] reg443 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg440 = (1'h0);
  reg [(5'h13):(1'h0)] reg439 = (1'h0);
  reg [(5'h12):(1'h0)] reg438 = (1'h0);
  reg [(4'h9):(1'h0)] reg437 = (1'h0);
  reg [(4'he):(1'h0)] reg435 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg434 = (1'h0);
  reg [(3'h4):(1'h0)] reg431 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar429 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg427 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar420 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar421 = (1'h0);
  reg [(3'h5):(1'h0)] reg420 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar417 = (1'h0);
  assign y = {wire469,
                 wire468,
                 wire416,
                 wire415,
                 reg467,
                 reg465,
                 reg463,
                 reg462,
                 reg458,
                 reg457,
                 reg455,
                 reg454,
                 reg452,
                 reg451,
                 reg450,
                 reg444,
                 reg442,
                 reg441,
                 reg436,
                 reg433,
                 reg432,
                 reg430,
                 reg428,
                 reg421,
                 reg426,
                 reg425,
                 reg424,
                 reg423,
                 reg422,
                 reg419,
                 reg418,
                 reg466,
                 reg464,
                 reg461,
                 reg460,
                 reg459,
                 reg456,
                 reg453,
                 forvar449,
                 reg448,
                 reg447,
                 reg446,
                 reg445,
                 reg443,
                 reg440,
                 reg439,
                 reg438,
                 reg437,
                 reg435,
                 reg434,
                 reg431,
                 forvar429,
                 reg427,
                 forvar420,
                 forvar421,
                 reg420,
                 forvar417,
                 (1'h0)};
  assign wire415 = ((8'hb6) ?
                       (wire414 << $signed((((8'h9d) << wire411) ?
                           $unsigned(wire410) : $signed(wire411)))) : wire410);
  assign wire416 = ((-$unsigned($signed((!(8'hb8))))) ?
                       ({(|wire414[(3'h7):(1'h0)]),
                               $unsigned($unsigned(wire412))} ?
                           wire410 : ((wire410[(2'h2):(2'h2)] >> wire412) ^ (wire412[(4'ha):(4'h8)] ?
                               (8'ha1) : $signed((8'ha2))))) : wire412);
  always
    @(posedge clk) begin
      for (forvar417 = (1'h0); (forvar417 < (1'h0)); forvar417 = (forvar417 + (1'h1)))
        begin
          if (wire410)
            begin
              reg418 <= $unsigned(($signed($signed((|wire410))) ?
                  wire416[(3'h5):(1'h0)] : (({wire410} ?
                          (8'ha6) : $unsigned(wire415)) ?
                      (wire410[(1'h0):(1'h0)] ?
                          $signed((8'ha4)) : wire411) : $signed({wire413}))));
              reg419 <= $unsigned($signed({wire416[(5'h13):(2'h2)]}));
            end
          else
            begin
              reg418 <= $signed(((-(-(reg418 && reg419))) <<< $unsigned($signed($unsigned((8'h9d))))));
            end
        end
      if ((~^(~^$unsigned(wire412))))
        begin
          reg420 = (!"B8po65EhON7U4hKXF0an");
          for (forvar421 = (1'h0); (forvar421 < (3'h4)); forvar421 = (forvar421 + (1'h1)))
            begin
              reg422 <= $signed({((wire416 && (wire412 ? (8'h9e) : (8'ha1))) ?
                      (^(forvar421 ?
                          wire415 : wire413)) : $unsigned($unsigned(wire413)))});
              reg423 <= $unsigned($unsigned(((wire414 ?
                  wire412[(4'ha):(2'h2)] : (wire415 ?
                      reg420 : wire410)) ~^ {(~&reg419)})));
              reg424 <= {((8'h9f) ?
                      (~^(|$signed(wire411))) : (({reg418,
                          wire414} <<< (+(8'ha5))) ^ $signed(wire411)))};
              reg425 <= (+(~&$unsigned(reg420[(1'h0):(1'h0)])));
              reg426 <= ((~^{($signed(wire416) ? $unsigned((8'haa)) : (8'ha4)),
                  $signed(reg420[(2'h3):(1'h0)])}) >= (~&reg425[(1'h1):(1'h1)]));
            end
        end
      else
        begin
          for (forvar420 = (1'h0); (forvar420 < (3'h4)); forvar420 = (forvar420 + (1'h1)))
            begin
              reg421 <= reg419[(4'he):(3'h6)];
              reg422 <= ($unsigned({($signed(reg426) == (~|wire414))}) & $signed($unsigned((8'hbc))));
              reg427 = $signed((reg422[(4'h8):(3'h5)] > wire411[(3'h4):(2'h3)]));
              reg428 <= (-((forvar421 == ($unsigned(wire411) < (~wire414))) ?
                  ((((8'ha2) & wire415) - (wire416 & (8'h9f))) ?
                      reg420 : reg418[(4'h8):(3'h6)]) : $signed($unsigned(wire413))));
            end
          for (forvar429 = (1'h0); (forvar429 < (2'h2)); forvar429 = (forvar429 + (1'h1)))
            begin
              reg430 <= ((reg419[(4'h8):(2'h2)] ?
                      reg422[(4'hc):(1'h1)] : $signed(((wire415 >= wire415) * {forvar420,
                          reg427}))) ?
                  reg426[(3'h6):(3'h4)] : (reg418 ?
                      wire410 : (^~$unsigned((reg424 ~^ wire414)))));
              reg431 = $unsigned((&wire412[(4'h8):(3'h5)]));
              reg432 <= (8'hba);
              reg433 <= $unsigned(($unsigned(((~(8'hbf)) ?
                      (reg424 >>> forvar420) : (&reg431))) ?
                  ($unsigned((~&reg418)) + (^~(reg427 ?
                      forvar417 : forvar417))) : {(&forvar417[(3'h5):(2'h3)])}));
            end
          if (($signed("VOTi6P4Px1JMQcu") & (+$signed("zP1RQMT3"))))
            begin
              reg434 = {((wire412 ?
                      $unsigned($signed((8'hb2))) : (+"PMe8DxFvMGGv6Fou")) >>> "H1wF1"),
                  $unsigned(forvar420)};
              reg435 = reg431;
              reg436 <= {(reg428 + reg428[(5'h10):(4'ha)])};
              reg437 = $signed(reg424);
              reg438 = wire416[(5'h13):(3'h6)];
            end
          else
            begin
              reg436 <= ($unsigned($signed((wire414 == reg426[(3'h6):(3'h4)]))) * reg426[(1'h0):(1'h0)]);
            end
          if (((reg435 ?
              (reg435 ~^ $signed($unsigned((8'haa)))) : $unsigned(reg438[(4'hc):(4'h8)])) == $unsigned($signed(reg432[(3'h6):(3'h6)]))))
            begin
              reg439 = ($unsigned((+$unsigned(reg419[(1'h1):(1'h0)]))) ?
                  {reg431[(1'h1):(1'h1)]} : (forvar421 ?
                      ((reg436 <= (reg431 >>> (8'haa))) ?
                          $unsigned((^wire413)) : (~&wire412)) : "KYL1ODL0krYeTId"));
              reg440 = reg435;
              reg441 <= $unsigned(((wire416[(3'h7):(1'h1)] ?
                      "07rV47CQr" : {reg419}) ?
                  wire416 : "dvZal"));
              reg442 <= $unsigned((^~((reg437 ?
                      forvar429[(4'ha):(4'h8)] : $signed((8'ha5))) ?
                  {reg431} : ((~reg424) ? reg439 : $unsigned((8'hbe))))));
            end
          else
            begin
              reg441 <= (forvar420 && (!(~^{reg437[(2'h3):(2'h3)]})));
              reg443 = $signed($unsigned((~$signed(reg434[(2'h2):(1'h0)]))));
              reg444 <= reg418;
              reg445 = forvar429;
              reg446 = reg443[(2'h3):(1'h1)];
            end
          reg447 = (((((~reg422) ?
                  forvar417 : (wire412 & reg422)) == (~|$signed(wire414))) ?
              (~&(-reg420)) : {({reg418} ? {forvar421} : $unsigned(forvar417)),
                  reg423}) >= (|({reg433[(3'h6):(1'h1)]} ?
              $signed({(8'ha3)}) : reg423[(3'h4):(2'h3)])));
        end
      reg448 = ($unsigned(reg442[(3'h4):(2'h3)]) ?
          $signed(($unsigned((8'ha1)) << $unsigned((reg420 ?
              (8'hac) : wire412)))) : reg446);
    end
  always
    @(posedge clk) begin
      for (forvar449 = (1'h0); (forvar449 < (2'h3)); forvar449 = (forvar449 + (1'h1)))
        begin
          reg450 <= $signed(reg441[(3'h5):(1'h1)]);
          reg451 <= $unsigned((8'h9e));
          reg452 <= (wire416 - "WdHabSiRQtDhI");
          reg453 = (~^$unsigned(($signed(reg426) > $unsigned((reg421 | reg430)))));
          if (reg418)
            begin
              reg454 <= {$unsigned((-wire415)),
                  ($signed((~&((8'hb8) ?
                      (8'hb3) : reg419))) + $unsigned(reg418))};
              reg455 <= ((~{{reg450, (reg421 ? reg423 : wire416)},
                  $unsigned($unsigned(reg452))}) >>> ((-wire414) ?
                  (|($signed(reg428) <<< (reg430 && reg430))) : ((+(~^reg453)) ?
                      ($signed(wire413) ?
                          wire411 : (reg451 ?
                              reg454 : reg428)) : ($unsigned(reg419) ?
                          (^reg444) : (wire412 ? wire413 : wire410)))));
              reg456 = wire413[(1'h0):(1'h0)];
            end
          else
            begin
              reg456 = (($unsigned(((reg442 != wire415) & (~|reg456))) != reg432) == $signed(((8'hba) >> reg422[(4'h9):(3'h7)])));
              reg457 <= reg432[(3'h6):(3'h5)];
              reg458 <= $unsigned((reg432 ?
                  $unsigned(reg453) : $signed($unsigned((reg425 >> wire410)))));
              reg459 = (reg436 >>> (^$unsigned((8'hb2))));
              reg460 = reg450[(3'h4):(3'h4)];
            end
        end
      if ($signed({$signed(reg456[(1'h0):(1'h0)])}))
        begin
          reg461 = {$unsigned(wire413[(4'hd):(4'hc)])};
          if ($unsigned(($unsigned(($signed(wire414) - reg423)) + reg432[(4'hb):(4'h9)])))
            begin
              reg462 <= reg422;
              reg463 <= (+(~|(((reg423 >> reg456) ?
                  (8'hae) : reg450) <<< reg432[(2'h3):(2'h2)])));
            end
          else
            begin
              reg464 = ({"sIsaaBuv6ePX6IZ",
                  ($unsigned((reg452 + (8'hba))) || (8'h9c))} <= $signed((reg456[(3'h6):(2'h3)] | ((~|reg442) ?
                  $unsigned(reg463) : (reg426 >> wire414)))));
            end
          reg465 <= ($signed(reg424[(2'h3):(1'h0)]) <<< (8'h9c));
        end
      else
        begin
          if ({((8'hb7) ?
                  $unsigned($unsigned((wire412 ?
                      reg426 : wire411))) : ((~^{(8'hb3)}) >= ((wire414 ?
                      (8'hbc) : (8'ha4)) && $unsigned(reg459))))})
            begin
              reg462 <= $unsigned($signed(reg423));
              reg463 <= {reg456[(3'h6):(2'h2)]};
              reg465 <= {(-($unsigned((|wire414)) <<< reg458))};
            end
          else
            begin
              reg461 = wire416[(4'hc):(4'h9)];
              reg462 <= reg463;
              reg464 = reg422;
              reg466 = ("rHlmHmbVKuzEMA6xEncV" ~^ reg424[(1'h1):(1'h1)]);
            end
          reg467 <= $signed($unsigned($unsigned((~&$unsigned(wire415)))));
        end
    end
  assign wire468 = wire416;
  assign wire469 = reg450;
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module275
#(parameter param384 = (~&(({{(8'h9c), (8'ha5)}} || (((8'ha5) ? (8'h9f) : (8'ha3)) > {(8'hb4)})) ? (|((&(8'hb3)) ^ ((8'hb7) ^~ (8'h9f)))) : (&({(8'haf)} ? (~|(8'hae)) : (~|(8'hbf)))))))
(y, clk, wire280, wire279, wire278, wire277, wire276);
  output wire [(32'h4ef):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire280;
  input wire [(4'hc):(1'h0)] wire279;
  input wire [(4'hf):(1'h0)] wire278;
  input wire signed [(5'h11):(1'h0)] wire277;
  input wire signed [(3'h4):(1'h0)] wire276;
  wire signed [(4'hd):(1'h0)] wire383;
  wire signed [(4'hf):(1'h0)] wire382;
  wire [(4'hd):(1'h0)] wire381;
  wire [(4'hd):(1'h0)] wire379;
  wire [(2'h2):(1'h0)] wire378;
  wire signed [(4'hc):(1'h0)] wire281;
  reg signed [(5'h10):(1'h0)] reg377 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg376 = (1'h0);
  reg [(4'hc):(1'h0)] reg375 = (1'h0);
  reg [(4'he):(1'h0)] reg367 = (1'h0);
  reg [(3'h5):(1'h0)] reg372 = (1'h0);
  reg [(3'h7):(1'h0)] reg370 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg369 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg365 = (1'h0);
  reg [(4'hb):(1'h0)] reg364 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg358 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg357 = (1'h0);
  reg [(3'h5):(1'h0)] reg355 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg349 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg348 = (1'h0);
  reg [(4'h9):(1'h0)] reg346 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg345 = (1'h0);
  reg [(3'h4):(1'h0)] reg344 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg343 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg338 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg337 = (1'h0);
  reg [(5'h11):(1'h0)] reg335 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg334 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg333 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg332 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg330 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg327 = (1'h0);
  reg signed [(4'he):(1'h0)] reg326 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg325 = (1'h0);
  reg [(4'he):(1'h0)] reg324 = (1'h0);
  reg [(2'h2):(1'h0)] reg323 = (1'h0);
  reg [(4'hd):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg319 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg316 = (1'h0);
  reg [(5'h11):(1'h0)] reg315 = (1'h0);
  reg [(5'h12):(1'h0)] reg313 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg311 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg305 = (1'h0);
  reg [(4'ha):(1'h0)] reg304 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg303 = (1'h0);
  reg [(4'he):(1'h0)] reg302 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg301 = (1'h0);
  reg [(5'h14):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg298 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg295 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg292 = (1'h0);
  reg signed [(4'he):(1'h0)] reg290 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg289 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg286 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg380 = (1'h0);
  reg [(2'h3):(1'h0)] forvar374 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar373 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg371 = (1'h0);
  reg [(4'hf):(1'h0)] reg368 = (1'h0);
  reg [(4'he):(1'h0)] forvar367 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg366 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg363 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar362 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg361 = (1'h0);
  reg [(4'hf):(1'h0)] reg360 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg359 = (1'h0);
  reg [(4'ha):(1'h0)] reg356 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar354 = (1'h0);
  reg [(4'hb):(1'h0)] reg353 = (1'h0);
  reg [(2'h2):(1'h0)] reg352 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg351 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg350 = (1'h0);
  reg [(5'h11):(1'h0)] forvar347 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar342 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg340 = (1'h0);
  reg [(3'h5):(1'h0)] forvar339 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg336 = (1'h0);
  reg signed [(4'he):(1'h0)] reg331 = (1'h0);
  reg [(5'h12):(1'h0)] reg329 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar328 = (1'h0);
  reg [(5'h11):(1'h0)] forvar321 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar320 = (1'h0);
  reg [(5'h12):(1'h0)] reg318 = (1'h0);
  reg [(5'h10):(1'h0)] reg317 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg314 = (1'h0);
  reg [(4'h9):(1'h0)] reg310 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg309 = (1'h0);
  reg [(4'h8):(1'h0)] reg308 = (1'h0);
  reg [(5'h15):(1'h0)] forvar307 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar306 = (1'h0);
  reg [(4'hd):(1'h0)] reg299 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg297 = (1'h0);
  reg [(5'h14):(1'h0)] forvar296 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg294 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar293 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg291 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar287 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg288 = (1'h0);
  reg [(4'hf):(1'h0)] reg285 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg284 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg283 = (1'h0);
  reg [(4'h9):(1'h0)] forvar282 = (1'h0);
  assign y = {wire383,
                 wire382,
                 wire381,
                 wire379,
                 wire378,
                 wire281,
                 reg377,
                 reg376,
                 reg375,
                 reg367,
                 reg372,
                 reg370,
                 reg369,
                 reg365,
                 reg364,
                 reg358,
                 reg357,
                 reg355,
                 reg349,
                 reg348,
                 reg346,
                 reg345,
                 reg344,
                 reg343,
                 reg341,
                 reg338,
                 reg337,
                 reg335,
                 reg334,
                 reg333,
                 reg332,
                 reg330,
                 reg327,
                 reg326,
                 reg325,
                 reg324,
                 reg323,
                 reg322,
                 reg319,
                 reg316,
                 reg315,
                 reg313,
                 reg312,
                 reg311,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg298,
                 reg295,
                 reg292,
                 reg290,
                 reg289,
                 reg287,
                 reg286,
                 reg380,
                 forvar374,
                 forvar373,
                 reg371,
                 reg368,
                 forvar367,
                 reg366,
                 reg363,
                 forvar362,
                 reg361,
                 reg360,
                 reg359,
                 reg356,
                 forvar354,
                 reg353,
                 reg352,
                 reg351,
                 reg350,
                 forvar347,
                 forvar342,
                 reg340,
                 forvar339,
                 reg336,
                 reg331,
                 reg329,
                 forvar328,
                 forvar321,
                 forvar320,
                 reg318,
                 reg317,
                 reg314,
                 reg310,
                 reg309,
                 reg308,
                 forvar307,
                 forvar306,
                 reg299,
                 reg297,
                 forvar296,
                 reg294,
                 forvar293,
                 reg291,
                 forvar287,
                 reg288,
                 reg285,
                 reg284,
                 reg283,
                 forvar282,
                 (1'h0)};
  assign wire281 = {$signed((((wire280 ?
                               wire279 : wire280) & $signed(wire276)) ?
                           $unsigned((-wire277)) : "Vx4dQDkzvQu4"))};
  always
    @(posedge clk) begin
      if (wire279[(4'hb):(3'h4)])
        begin
          for (forvar282 = (1'h0); (forvar282 < (1'h0)); forvar282 = (forvar282 + (1'h1)))
            begin
              reg283 = wire277;
              reg284 = wire276[(3'h4):(3'h4)];
            end
          if (($signed($signed(forvar282)) ?
              (&$signed(wire276[(2'h3):(1'h1)])) : (forvar282 << wire281)))
            begin
              reg285 = wire278;
              reg286 <= reg285[(1'h1):(1'h0)];
              reg287 <= (~^$signed(($unsigned((wire280 >> wire278)) ?
                  ("mFIagbFy" + ((8'ha6) * wire279)) : "1IhJa64KovINnrfQUq")));
            end
          else
            begin
              reg285 = $unsigned($unsigned($unsigned(wire277)));
              reg286 <= $unsigned(wire280[(4'ha):(2'h2)]);
              reg287 <= $signed($signed((^(wire279[(3'h7):(2'h2)] <<< wire280[(4'hf):(4'he)]))));
              reg288 = $signed(wire277);
              reg289 <= $unsigned(({(8'hbe)} ?
                  (((~&reg288) ? reg286 : wire278) ?
                      reg283 : {$signed(reg286)}) : wire276[(2'h2):(2'h2)]));
            end
        end
      else
        begin
          for (forvar282 = (1'h0); (forvar282 < (2'h2)); forvar282 = (forvar282 + (1'h1)))
            begin
              reg286 <= reg286[(5'h10):(4'h9)];
            end
          for (forvar287 = (1'h0); (forvar287 < (2'h2)); forvar287 = (forvar287 + (1'h1)))
            begin
              reg288 = $unsigned($unsigned(reg283[(4'hf):(4'hb)]));
              reg289 <= ({$signed((reg287[(3'h4):(2'h2)] ?
                      $unsigned(reg288) : (reg289 | reg284))),
                  $unsigned(reg286[(2'h2):(1'h1)])} > {(((wire281 ?
                              (8'ha6) : forvar282) ?
                          "UWXo1T" : (-(8'hb7))) ?
                      $signed((reg289 <= wire278)) : {{(8'hb7)}})});
              reg290 <= $signed($signed(wire281));
            end
          reg291 = wire277[(4'hf):(1'h1)];
          reg292 <= $unsigned(wire277);
        end
      for (forvar293 = (1'h0); (forvar293 < (2'h3)); forvar293 = (forvar293 + (1'h1)))
        begin
          reg294 = forvar293;
          reg295 <= $signed((&(((8'hb1) ?
                  wire279[(4'hc):(3'h5)] : reg284[(3'h5):(1'h1)]) ?
              (reg290[(1'h1):(1'h1)] ?
                  reg291[(4'hc):(3'h4)] : forvar282[(3'h4):(1'h1)]) : $signed({wire281,
                  (8'ha0)}))));
          for (forvar296 = (1'h0); (forvar296 < (1'h0)); forvar296 = (forvar296 + (1'h1)))
            begin
              reg297 = (((reg287 ?
                          forvar287 : ((+reg292) <<< (forvar287 ?
                              (8'hb5) : reg289))) ?
                      reg295 : reg292[(4'h9):(2'h2)]) ?
                  "0WTDX8J" : ({{(forvar282 + wire278), $signed(reg291)}} ?
                      reg285[(3'h4):(2'h2)] : wire280[(4'hf):(3'h7)]));
              reg298 <= wire278[(1'h1):(1'h1)];
              reg299 = $unsigned($signed(reg292));
              reg300 <= ((!($unsigned((^(8'hb0))) ?
                      ($signed(wire280) ?
                          ((7'h41) ?
                              wire280 : reg285) : $unsigned(reg284)) : $unsigned(reg286[(4'he):(3'h4)]))) ?
                  (((~^(&reg290)) ?
                      (8'ha9) : (~|reg283[(1'h0):(1'h0)])) >>> wire281[(4'ha):(4'h9)]) : reg285[(4'hf):(4'hf)]);
            end
          if ($unsigned(reg283))
            begin
              reg301 <= "qMSL";
              reg302 <= (^(~^wire276));
              reg303 <= $unsigned(reg295[(3'h7):(1'h0)]);
              reg304 <= (^~({(reg299[(4'ha):(3'h7)] ?
                      (~reg291) : reg292[(1'h1):(1'h0)])} | (~^(~&(~&(8'ha5))))));
              reg305 <= reg284;
            end
          else
            begin
              reg301 <= $unsigned({(((reg289 ?
                      wire279 : reg284) | $unsigned(reg288)) >>> ((&wire280) || (-reg291)))});
            end
        end
      for (forvar306 = (1'h0); (forvar306 < (1'h0)); forvar306 = (forvar306 + (1'h1)))
        begin
          for (forvar307 = (1'h0); (forvar307 < (1'h0)); forvar307 = (forvar307 + (1'h1)))
            begin
              reg308 = forvar306[(4'hc):(3'h5)];
              reg309 = $signed(($unsigned(reg288) ?
                  $signed($signed({wire280})) : ("nzSWkYGvxa" ?
                      "7iX2irqHRN99grMn" : $unsigned(reg301))));
            end
          reg310 = reg299[(1'h0):(1'h0)];
          if ((&(|{forvar296[(1'h0):(1'h0)],
              ($unsigned(reg291) || $unsigned(wire280))})))
            begin
              reg311 <= ((|(~^(~^reg298))) && (^~$signed((reg295[(3'h7):(1'h1)] ?
                  (wire279 ? reg288 : reg291) : reg303[(1'h0):(1'h0)]))));
              reg312 <= wire281[(4'hb):(4'h8)];
              reg313 <= (^reg311);
            end
          else
            begin
              reg311 <= ((|((reg304[(3'h5):(3'h4)] < $signed(reg298)) ?
                      {reg290,
                          reg285[(4'hd):(3'h6)]} : (forvar293[(1'h0):(1'h0)] >= (reg304 & forvar307)))) ?
                  (-($unsigned($signed(reg313)) & (8'haf))) : reg301);
              reg314 = forvar293;
              reg315 <= ({forvar293[(2'h3):(2'h2)]} != reg308[(2'h2):(1'h0)]);
              reg316 <= ($signed(((reg301 ?
                      $signed(reg283) : wire281[(4'ha):(2'h2)]) - ((~reg304) ?
                      (&reg313) : (|reg309)))) ?
                  $unsigned(((~((8'hbb) >= (8'ha7))) ?
                      ((reg288 ?
                          reg314 : reg309) - $signed((8'ha4))) : "oFRZgw")) : ($unsigned(reg294[(5'h10):(3'h7)]) ?
                      reg302 : (($signed(reg298) ? reg288 : reg291) ?
                          $signed($unsigned(reg290)) : $signed((~reg303)))));
              reg317 = ($unsigned({wire277[(4'h9):(1'h0)]}) >> $signed((reg295[(3'h7):(3'h5)] ?
                  {{wire280},
                      wire276[(2'h2):(2'h2)]} : (forvar293[(2'h2):(1'h1)] ?
                      ((8'hbc) + reg288) : {reg300, reg315}))));
            end
          reg318 = (~^$unsigned($unsigned(reg286[(4'h8):(3'h4)])));
        end
    end
  always
    @(posedge clk) begin
      reg319 <= ($unsigned({$unsigned({(8'hbd), reg287}),
              ({reg298, wire277} <<< wire278[(3'h5):(1'h1)])}) ?
          (|reg301[(5'h10):(4'hb)]) : $unsigned((~reg316[(5'h12):(1'h0)])));
      for (forvar320 = (1'h0); (forvar320 < (1'h1)); forvar320 = (forvar320 + (1'h1)))
        begin
          for (forvar321 = (1'h0); (forvar321 < (1'h1)); forvar321 = (forvar321 + (1'h1)))
            begin
              reg322 <= (~|$unsigned((8'hb6)));
              reg323 <= $unsigned(reg290[(4'h8):(3'h4)]);
              reg324 <= {(reg315 <= wire281[(4'h9):(2'h2)])};
            end
          reg325 <= reg319[(1'h1):(1'h1)];
          if ((~reg322[(3'h7):(1'h1)]))
            begin
              reg326 <= (reg292 ?
                  (reg292[(4'h8):(1'h0)] * ($signed(wire280) ?
                      reg301 : (!$signed(wire279)))) : (~^$unsigned($signed((reg298 ?
                      reg322 : reg311)))));
              reg327 <= (forvar321 <= $unsigned(($signed((^~wire278)) ?
                  wire276[(1'h0):(1'h0)] : $signed($signed(reg315)))));
            end
          else
            begin
              reg326 <= reg303;
            end
          for (forvar328 = (1'h0); (forvar328 < (1'h1)); forvar328 = (forvar328 + (1'h1)))
            begin
              reg329 = $signed((!($signed(((8'haa) * reg303)) ?
                  (reg319 ? $unsigned(reg292) : (&(7'h43))) : (~|(8'hb9)))));
              reg330 <= $signed((reg287 ^ ($signed($unsigned(wire278)) <= (wire277 - reg290))));
              reg331 = $unsigned(wire276);
              reg332 <= $unsigned(wire277);
            end
        end
      if ((reg290 + reg311[(1'h0):(1'h0)]))
        begin
          reg333 <= $unsigned((reg324 ? reg326 : reg290[(4'h9):(3'h6)]));
          reg334 <= (^~$unsigned($signed($signed(reg301[(5'h12):(5'h11)]))));
          reg335 <= (+($unsigned($signed((^reg290))) ?
              {"WLqYxnR3Ql"} : reg333));
        end
      else
        begin
          reg333 <= $unsigned(reg305);
          if ($signed(wire280[(4'hf):(2'h2)]))
            begin
              reg336 = ((reg325 ?
                      (~|((reg315 ^ (8'hab)) ?
                          "76qDZAGJrD" : ((8'hb1) >= forvar320))) : $unsigned(reg300[(4'hf):(4'h9)])) ?
                  reg301[(4'hf):(3'h4)] : ((({reg319} >> reg329) | ($signed(reg326) == (-(8'ha7)))) ?
                      (((reg289 ? reg315 : reg312) ?
                          {reg319,
                              reg332} : (forvar321 || reg329)) ^~ (wire276[(3'h4):(1'h1)] >>> $unsigned(reg286))) : "IaBGX7XaIn"));
              reg337 <= reg322;
            end
          else
            begin
              reg334 <= (|{({(reg289 ^ reg333)} ~^ ($unsigned((8'hbf)) ?
                      $unsigned((8'ha7)) : "C8bOk2NBdxMi9"))});
            end
          reg338 <= wire277;
          for (forvar339 = (1'h0); (forvar339 < (2'h2)); forvar339 = (forvar339 + (1'h1)))
            begin
              reg340 = $unsigned(wire276);
              reg341 <= "KLfkQ7MAiWMV";
            end
          for (forvar342 = (1'h0); (forvar342 < (1'h1)); forvar342 = (forvar342 + (1'h1)))
            begin
              reg343 <= (wire279 ?
                  ((($unsigned(reg289) ? reg312[(5'h10):(4'hc)] : {reg319}) ?
                      reg337 : $unsigned(reg300)) ^~ $signed(((forvar342 - reg338) | (reg340 ?
                      reg327 : reg286)))) : forvar328[(4'h8):(1'h0)]);
              reg344 <= $unsigned((7'h44));
              reg345 <= $signed((~{(^(&reg289))}));
              reg346 <= wire281;
            end
        end
      for (forvar347 = (1'h0); (forvar347 < (3'h4)); forvar347 = (forvar347 + (1'h1)))
        begin
          reg348 <= $signed(wire279[(3'h6):(1'h1)]);
          if ($signed($unsigned($signed({"5a9hH7Uvna8fp2Ylbw",
              (reg326 ? reg304 : reg338)}))))
            begin
              reg349 <= ($unsigned(((wire278 >>> $signed(reg316)) >> wire279[(4'h8):(4'h8)])) ?
                  (!($signed("M0rsbdYHV1uA1UvVf2") ~^ ($signed(reg340) ?
                      (~^wire276) : reg332[(1'h1):(1'h0)]))) : reg319);
              reg350 = reg319[(1'h0):(1'h0)];
              reg351 = $unsigned(((reg343[(4'hd):(4'h9)] || ((reg319 ?
                      reg331 : reg350) << reg295[(4'ha):(4'ha)])) ?
                  (8'hb9) : {{{(8'hbf)}, (reg329 ~^ (8'hbc))}}));
              reg352 = reg327[(2'h2):(1'h1)];
            end
          else
            begin
              reg350 = reg312;
            end
          reg353 = ((wire280 ?
                  $unsigned(({reg345} + {reg287})) : ($signed(((8'hb3) && reg313)) ?
                      {$unsigned(reg338),
                          $unsigned(forvar321)} : (!((8'h9e) != reg343)))) ?
              forvar328[(1'h1):(1'h1)] : (!reg332));
        end
      for (forvar354 = (1'h0); (forvar354 < (2'h3)); forvar354 = (forvar354 + (1'h1)))
        begin
          if ($signed(reg346))
            begin
              reg355 <= (((!(-(reg289 ? reg302 : reg312))) ?
                  reg352[(2'h2):(2'h2)] : {$signed((~reg350))}) >> (($signed({reg298,
                      reg312}) * ($unsigned((8'haa)) - {(8'hac)})) ?
                  (~|((reg304 ? reg301 : reg350) ?
                      (8'hb1) : (~&forvar339))) : reg311[(2'h3):(1'h1)]));
              reg356 = ("7sx9LtrIeSHpA" == $unsigned({(reg286 ^~ $unsigned(reg338)),
                  reg295}));
              reg357 <= forvar321[(4'hb):(1'h1)];
            end
          else
            begin
              reg355 <= ($signed($unsigned(((wire281 ?
                  (8'hbb) : reg348) <<< $unsigned(reg305)))) & ((8'h9f) ?
                  ((~^(&forvar320)) ?
                      "NiGNbCerCOmfgxGi5nhw" : forvar339[(3'h4):(3'h4)]) : reg356[(4'ha):(4'ha)]));
              reg357 <= $signed((!(($unsigned(reg326) >= $unsigned(reg302)) < reg344)));
              reg358 <= wire281[(3'h6):(3'h4)];
              reg359 = $unsigned({$signed($signed($unsigned(reg312))),
                  $unsigned(({forvar347, reg289} >= (wire280 != wire281)))});
            end
          reg360 = ((($signed((8'hbe)) && (reg351 >= (forvar328 + reg340))) >> (&wire278)) - (forvar354[(2'h2):(1'h1)] != reg327));
          reg361 = $signed({$unsigned($unsigned($signed(reg313))),
              {(|$unsigned(reg304)), (~^(reg359 ? reg326 : reg329))}});
          for (forvar362 = (1'h0); (forvar362 < (2'h3)); forvar362 = (forvar362 + (1'h1)))
            begin
              reg363 = (reg325 ?
                  ((!((reg316 ? reg302 : reg290) ?
                          reg312 : $unsigned(reg311))) ?
                      ($signed($signed(reg327)) ?
                          ((^reg290) ?
                              (~reg351) : (reg311 - reg322)) : $unsigned($unsigned(reg329))) : (8'hab)) : ($unsigned($signed((reg336 || reg345))) ?
                      $unsigned(((reg353 ? (8'hb2) : reg304) ?
                          {wire276} : $signed(reg345))) : $signed($signed((8'h9f)))));
              reg364 <= $unsigned(reg348);
              reg365 <= $signed((reg355 ~^ $signed((reg338 + wire276))));
              reg366 = (&(reg364 <= (reg363[(1'h0):(1'h0)] ?
                  reg334 : ((!reg335) ? {reg336, wire278} : {(8'hbe)}))));
            end
        end
    end
  always
    @(posedge clk) begin
      if ((reg311 ^~ reg327[(1'h1):(1'h0)]))
        begin
          for (forvar367 = (1'h0); (forvar367 < (2'h3)); forvar367 = (forvar367 + (1'h1)))
            begin
              reg368 = $signed((reg300 ?
                  {""} : (~&(~(reg302 ? wire280 : (8'haf))))));
              reg369 <= $unsigned(((~|({reg333} >= $signed(reg319))) ?
                  {((~wire278) ?
                          reg349 : (reg292 ^ (8'hb2)))} : reg290[(4'h8):(3'h6)]));
            end
          reg370 <= reg334[(5'h13):(4'hb)];
          reg371 = $unsigned((reg346[(4'h9):(4'h9)] ?
              {reg302[(2'h2):(2'h2)]} : $signed((((8'hb2) <= (8'ha1)) ?
                  {reg295, reg368} : $signed((8'h9f))))));
          reg372 <= reg338;
        end
      else
        begin
          reg367 <= reg286;
        end
      for (forvar373 = (1'h0); (forvar373 < (2'h2)); forvar373 = (forvar373 + (1'h1)))
        begin
          for (forvar374 = (1'h0); (forvar374 < (2'h3)); forvar374 = (forvar374 + (1'h1)))
            begin
              reg375 <= forvar373[(4'hd):(2'h3)];
              reg376 <= $signed(reg369);
            end
          reg377 <= reg367;
        end
    end
  assign wire378 = (reg370 < ((((reg333 ?
                       reg357 : reg327) ^ reg300) <= (^~reg377[(4'hf):(4'he)])) <= ($unsigned(reg295[(3'h6):(1'h1)]) ?
                       ($signed(reg322) ?
                           ((8'ha4) ? reg358 : reg301) : (8'had)) : ((reg292 ?
                               (8'ha1) : reg295) ?
                           $signed(reg301) : reg333[(4'hc):(4'hb)]))));
  assign wire379 = ($signed($unsigned((reg338[(5'h14):(2'h2)] >= $unsigned(reg292)))) ?
                       ((reg330[(2'h2):(2'h2)] >= (&$unsigned((8'ha0)))) ?
                           reg313[(3'h4):(3'h4)] : reg346[(2'h3):(2'h3)]) : ("rYqdfOb" ~^ reg326));
  always
    @(posedge clk) begin
      reg380 = reg311[(1'h1):(1'h1)];
    end
  assign wire381 = reg343[(4'hc):(1'h1)];
  assign wire382 = $unsigned(reg348);
  assign wire383 = (+{{$unsigned($unsigned(reg349))}, reg303});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module172  (y, clk, wire176, wire175, wire174, wire173);
  output wire [(32'h47c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire176;
  input wire [(3'h7):(1'h0)] wire175;
  input wire [(4'hc):(1'h0)] wire174;
  input wire signed [(3'h5):(1'h0)] wire173;
  wire [(4'h8):(1'h0)] wire213;
  wire [(2'h2):(1'h0)] wire212;
  wire [(4'h9):(1'h0)] wire201;
  wire [(5'h10):(1'h0)] wire200;
  wire signed [(4'he):(1'h0)] wire199;
  wire signed [(4'h9):(1'h0)] wire179;
  wire [(3'h6):(1'h0)] wire178;
  wire signed [(4'hd):(1'h0)] wire177;
  reg [(4'hf):(1'h0)] reg272 = (1'h0);
  reg [(4'hf):(1'h0)] reg271 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg270 = (1'h0);
  reg [(4'hf):(1'h0)] reg268 = (1'h0);
  reg [(4'hc):(1'h0)] reg267 = (1'h0);
  reg [(4'hd):(1'h0)] reg266 = (1'h0);
  reg [(2'h2):(1'h0)] reg265 = (1'h0);
  reg [(4'he):(1'h0)] reg264 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg262 = (1'h0);
  reg [(4'hb):(1'h0)] reg261 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg260 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg257 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg256 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg255 = (1'h0);
  reg signed [(4'he):(1'h0)] reg254 = (1'h0);
  reg [(4'h9):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg249 = (1'h0);
  reg [(5'h10):(1'h0)] reg248 = (1'h0);
  reg [(5'h14):(1'h0)] reg246 = (1'h0);
  reg [(4'hd):(1'h0)] reg244 = (1'h0);
  reg signed [(4'he):(1'h0)] reg243 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg240 = (1'h0);
  reg [(5'h15):(1'h0)] reg236 = (1'h0);
  reg [(5'h10):(1'h0)] reg235 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg233 = (1'h0);
  reg [(2'h3):(1'h0)] reg230 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg229 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg224 = (1'h0);
  reg [(4'ha):(1'h0)] reg223 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg219 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg218 = (1'h0);
  reg [(5'h15):(1'h0)] reg215 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg214 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg205 = (1'h0);
  reg [(5'h12):(1'h0)] reg209 = (1'h0);
  reg [(5'h14):(1'h0)] reg207 = (1'h0);
  reg [(4'hd):(1'h0)] reg204 = (1'h0);
  reg signed [(4'he):(1'h0)] reg202 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg198 = (1'h0);
  reg [(3'h7):(1'h0)] reg197 = (1'h0);
  reg [(5'h13):(1'h0)] reg196 = (1'h0);
  reg [(3'h6):(1'h0)] reg195 = (1'h0);
  reg [(3'h7):(1'h0)] reg191 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg192 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg190 = (1'h0);
  reg [(5'h13):(1'h0)] reg183 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg182 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg181 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg269 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg263 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg259 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar258 = (1'h0);
  reg [(4'hb):(1'h0)] reg247 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg253 = (1'h0);
  reg [(5'h14):(1'h0)] reg252 = (1'h0);
  reg [(3'h7):(1'h0)] reg251 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar247 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg245 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg242 = (1'h0);
  reg [(5'h14):(1'h0)] reg241 = (1'h0);
  reg [(4'ha):(1'h0)] forvar239 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg238 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg237 = (1'h0);
  reg [(2'h3):(1'h0)] forvar234 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar232 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar231 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg228 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg227 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar226 = (1'h0);
  reg [(5'h14):(1'h0)] reg225 = (1'h0);
  reg [(2'h2):(1'h0)] reg222 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg220 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar217 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar216 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg211 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg210 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar208 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg206 = (1'h0);
  reg [(4'he):(1'h0)] forvar205 = (1'h0);
  reg [(4'he):(1'h0)] reg203 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg194 = (1'h0);
  reg [(3'h5):(1'h0)] forvar193 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg187 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar191 = (1'h0);
  reg [(4'hf):(1'h0)] reg189 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg188 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar187 = (1'h0);
  reg [(3'h5):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg185 = (1'h0);
  reg [(4'hb):(1'h0)] reg184 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar180 = (1'h0);
  assign y = {wire213,
                 wire212,
                 wire201,
                 wire200,
                 wire199,
                 wire179,
                 wire178,
                 wire177,
                 reg272,
                 reg271,
                 reg270,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg264,
                 reg262,
                 reg261,
                 reg260,
                 reg257,
                 reg256,
                 reg255,
                 reg254,
                 reg250,
                 reg249,
                 reg248,
                 reg246,
                 reg244,
                 reg243,
                 reg240,
                 reg236,
                 reg235,
                 reg233,
                 reg230,
                 reg229,
                 reg224,
                 reg223,
                 reg219,
                 reg218,
                 reg215,
                 reg214,
                 reg205,
                 reg209,
                 reg207,
                 reg204,
                 reg202,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg191,
                 reg192,
                 reg190,
                 reg183,
                 reg182,
                 reg181,
                 reg269,
                 reg263,
                 reg259,
                 forvar258,
                 reg247,
                 reg253,
                 reg252,
                 reg251,
                 forvar247,
                 reg245,
                 reg242,
                 reg241,
                 forvar239,
                 reg238,
                 reg237,
                 forvar234,
                 forvar232,
                 forvar231,
                 reg228,
                 reg227,
                 forvar226,
                 reg225,
                 reg222,
                 reg221,
                 reg220,
                 forvar217,
                 forvar216,
                 reg208,
                 reg211,
                 reg210,
                 forvar208,
                 reg206,
                 forvar205,
                 reg203,
                 reg194,
                 forvar193,
                 reg187,
                 forvar191,
                 reg189,
                 reg188,
                 forvar187,
                 reg186,
                 reg185,
                 reg184,
                 forvar180,
                 (1'h0)};
  assign wire177 = ((~wire173) ?
                       $unsigned((~^({wire176} & $unsigned(wire176)))) : wire173[(2'h2):(1'h0)]);
  assign wire178 = {((^(((8'ha1) | wire175) ?
                               wire174[(1'h1):(1'h0)] : {wire177})) ?
                           $unsigned((&"LVSPwGAwG60xBA1")) : $signed($unsigned((wire174 ?
                               wire174 : wire177))))};
  assign wire179 = wire173[(2'h2):(1'h1)];
  always
    @(posedge clk) begin
      for (forvar180 = (1'h0); (forvar180 < (3'h4)); forvar180 = (forvar180 + (1'h1)))
        begin
          reg181 <= wire177;
        end
      if (wire175[(3'h4):(3'h4)])
        begin
          reg182 <= forvar180;
          reg183 <= wire178[(2'h2):(2'h2)];
        end
      else
        begin
          reg184 = "sJPLLY3ONd";
          reg185 = wire177;
        end
      reg186 = (wire176 != $signed(wire178));
      if (forvar180)
        begin
          for (forvar187 = (1'h0); (forvar187 < (1'h1)); forvar187 = (forvar187 + (1'h1)))
            begin
              reg188 = $signed((^~wire179[(3'h6):(2'h2)]));
            end
          reg189 = (+wire175[(1'h1):(1'h1)]);
          reg190 <= $unsigned(reg182[(1'h0):(1'h0)]);
          for (forvar191 = (1'h0); (forvar191 < (1'h1)); forvar191 = (forvar191 + (1'h1)))
            begin
              reg192 <= $signed($signed(wire176[(2'h2):(2'h2)]));
            end
        end
      else
        begin
          reg187 = ($signed(reg186) ?
              reg184 : (((8'hbb) && $unsigned(wire177[(3'h6):(1'h1)])) ?
                  ($signed({wire175,
                      wire173}) + (8'hb6)) : ((wire177[(1'h1):(1'h1)] ?
                          (reg181 >> (8'ha0)) : (wire174 ? reg185 : reg190)) ?
                      forvar191[(2'h2):(1'h1)] : (wire177 | $signed(wire177)))));
          reg190 <= (8'had);
          reg191 <= (&$signed((~|reg190[(1'h0):(1'h0)])));
        end
    end
  always
    @(posedge clk) begin
      for (forvar193 = (1'h0); (forvar193 < (2'h2)); forvar193 = (forvar193 + (1'h1)))
        begin
          if ((reg181 << wire179))
            begin
              reg194 = (reg190[(4'hd):(1'h1)] ?
                  reg192 : $signed($signed((8'ha7))));
              reg195 <= $signed(wire176[(2'h2):(1'h1)]);
              reg196 <= "DK";
            end
          else
            begin
              reg195 <= wire179[(4'h8):(4'h8)];
            end
        end
      reg197 <= $signed(({(reg190 && $signed((8'hb0)))} - wire176));
      reg198 <= ($signed($unsigned(wire176)) ?
          $unsigned(forvar193[(3'h5):(1'h1)]) : (wire175[(1'h1):(1'h0)] ?
              reg197 : (({reg181} && {reg192,
                  wire178}) >>> ((-wire177) & $unsigned(forvar193)))));
    end
  assign wire199 = $unsigned(reg192[(3'h6):(3'h4)]);
  assign wire200 = $signed($signed((wire179[(2'h2):(2'h2)] <= ($unsigned(reg195) > (reg191 ?
                       reg195 : (8'hb7))))));
  assign wire201 = {(wire178 ?
                           ($signed(wire199) ~^ $unsigned($unsigned(reg182))) : (~^wire177[(4'ha):(4'h9)]))};
  always
    @(posedge clk) begin
      reg202 <= {$unsigned(wire176[(1'h0):(1'h0)])};
      reg203 = $unsigned(wire177[(3'h7):(3'h6)]);
      reg204 <= (+wire179);
    end
  always
    @(posedge clk) begin
      if ((reg182[(1'h1):(1'h1)] - wire173))
        begin
          for (forvar205 = (1'h0); (forvar205 < (2'h3)); forvar205 = (forvar205 + (1'h1)))
            begin
              reg206 = (reg202 | (~^wire174));
              reg207 <= (({({reg204} >>> ((7'h40) ? wire177 : wire201)),
                  (8'hb8)} >> reg191[(3'h6):(2'h2)]) ~^ reg198[(3'h4):(1'h0)]);
            end
          for (forvar208 = (1'h0); (forvar208 < (1'h1)); forvar208 = (forvar208 + (1'h1)))
            begin
              reg209 <= (|"tLAL1hLYhh");
              reg210 = ({reg206[(3'h5):(2'h3)],
                      $unsigned((^$unsigned(forvar205)))} ?
                  $signed((8'ha6)) : ((reg196 <<< $signed((reg190 ?
                          (7'h40) : reg195))) ?
                      ((reg183 ? {(8'hae), reg209} : {reg206, (8'hb4)}) ?
                          $unsigned($unsigned(reg183)) : (reg190 != (wire177 ?
                              (8'hb4) : (8'hac)))) : reg204));
              reg211 = (((~|wire175[(1'h0):(1'h0)]) >> forvar208) != (|reg202[(1'h0):(1'h0)]));
            end
        end
      else
        begin
          if ({($signed((|(reg197 < wire200))) < {((forvar205 ?
                      reg190 : reg191) || (~&wire174))})})
            begin
              reg205 <= (wire179 <<< $signed($unsigned($signed((forvar205 <= reg204)))));
            end
          else
            begin
              reg206 = (forvar208 ?
                  (^~(((~&forvar208) >> (reg198 != reg209)) ?
                      {(^~(8'ha9)),
                          (8'hae)} : (^~$unsigned((7'h44))))) : forvar208[(1'h0):(1'h0)]);
              reg208 = $signed(wire199[(1'h1):(1'h1)]);
            end
        end
    end
  assign wire212 = (~&reg190);
  assign wire213 = ((wire200[(2'h3):(1'h0)] ?
                           $signed($unsigned((~&wire175))) : $signed("PR0EfXVrX")) ?
                       $signed(reg196[(3'h6):(1'h1)]) : "AixSxEBcFAh");
  always
    @(posedge clk) begin
      reg214 <= {(&(&reg207[(4'ha):(4'ha)]))};
      reg215 <= reg214;
      for (forvar216 = (1'h0); (forvar216 < (2'h2)); forvar216 = (forvar216 + (1'h1)))
        begin
          for (forvar217 = (1'h0); (forvar217 < (1'h0)); forvar217 = (forvar217 + (1'h1)))
            begin
              reg218 <= $unsigned($unsigned(wire175));
              reg219 <= (~reg202[(2'h2):(1'h1)]);
              reg220 = (^($signed(reg219[(1'h0):(1'h0)]) ?
                  $unsigned((reg204 ?
                      (wire175 ?
                          reg214 : reg181) : $unsigned(reg183))) : (~^(~|(wire199 ?
                      wire173 : wire173)))));
              reg221 = (^wire177[(4'hb):(4'h8)]);
              reg222 = $signed((reg204[(3'h4):(3'h4)] && wire174[(1'h1):(1'h0)]));
            end
          if ($unsigned($unsigned(((-wire175) == (~^$unsigned(reg197))))))
            begin
              reg223 <= ((((^~(reg214 - wire174)) == {(7'h44),
                          reg218[(4'ha):(3'h7)]}) ?
                      ((((7'h42) ? reg190 : wire213) ?
                          $signed(reg191) : $unsigned((7'h40))) == (&(wire213 ?
                          reg183 : wire200))) : $signed((7'h43))) ?
                  ($unsigned(reg221) ?
                      wire200 : reg205[(4'h9):(1'h1)]) : ($unsigned((8'ha4)) ?
                      ($unsigned(wire212) ?
                          wire199[(4'h8):(3'h4)] : ($unsigned(reg183) <<< "5Xzyioyfccg")) : reg218[(4'hc):(1'h0)]));
              reg224 <= $signed($signed(reg209));
              reg225 = $unsigned((reg224 * $unsigned($signed(reg223[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg223 <= reg222[(1'h1):(1'h0)];
              reg224 <= reg220[(3'h5):(1'h1)];
              reg225 = reg182;
            end
        end
      for (forvar226 = (1'h0); (forvar226 < (2'h2)); forvar226 = (forvar226 + (1'h1)))
        begin
          reg227 = reg195;
          reg228 = (^(+reg181[(3'h4):(1'h1)]));
          reg229 <= {(reg218[(4'ha):(3'h6)] ?
                  wire173 : $signed($signed((~^wire200)))),
              $unsigned((~^({reg207, forvar217} | $unsigned(reg183))))};
        end
      reg230 <= reg181[(2'h3):(2'h2)];
    end
  always
    @(posedge clk) begin
      for (forvar231 = (1'h0); (forvar231 < (1'h0)); forvar231 = (forvar231 + (1'h1)))
        begin
          for (forvar232 = (1'h0); (forvar232 < (2'h3)); forvar232 = (forvar232 + (1'h1)))
            begin
              reg233 <= (reg207 ? wire199[(4'hc):(4'ha)] : (8'ha1));
            end
          for (forvar234 = (1'h0); (forvar234 < (1'h0)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 <= wire200;
              reg236 <= (-reg230[(1'h0):(1'h0)]);
              reg237 = {$signed(reg235)};
            end
          reg238 = $unsigned((reg192 && (~|{(reg230 ? forvar232 : wire174)})));
          for (forvar239 = (1'h0); (forvar239 < (1'h0)); forvar239 = (forvar239 + (1'h1)))
            begin
              reg240 <= $unsigned(("" ?
                  wire199 : $signed(((^reg237) ?
                      $unsigned(reg205) : ((8'hb7) ? wire174 : reg191)))));
              reg241 = (wire173 >= (wire173[(3'h4):(1'h1)] ?
                  (8'ha5) : ($unsigned($signed((8'ha0))) ?
                      (reg233 >= $unsigned(wire173)) : wire179[(2'h3):(2'h2)])));
              reg242 = "kMKqCoFA";
              reg243 <= (reg190[(4'hf):(3'h7)] ?
                  (~|$unsigned(reg219[(3'h4):(1'h0)])) : reg229[(1'h0):(1'h0)]);
            end
          reg244 <= $signed($signed(((^~"c7AJzJHys2qF0") > ((wire177 >>> forvar232) ?
              $signed(reg218) : reg198[(3'h6):(1'h0)]))));
        end
      reg245 = forvar239[(3'h7):(3'h5)];
      if (($unsigned(({{reg202}} ?
              wire179[(2'h2):(2'h2)] : (|((8'hb7) ^~ forvar234)))) ?
          reg238 : reg183))
        begin
          reg246 <= $unsigned(reg215);
          for (forvar247 = (1'h0); (forvar247 < (2'h2)); forvar247 = (forvar247 + (1'h1)))
            begin
              reg248 <= forvar232;
              reg249 <= $signed(wire179);
              reg250 <= ($unsigned((|$unsigned(forvar231[(3'h5):(3'h4)]))) ^ {{((~^reg230) || (~wire200)),
                      (-reg238)}});
            end
          if ((~(((^~reg250) ?
              "kEN0a0awi4QgroE" : $signed($unsigned(reg192))) + {reg238})))
            begin
              reg251 = $unsigned(wire176);
              reg252 = (wire176[(1'h1):(1'h0)] ?
                  $signed(wire173) : $signed((8'ha3)));
              reg253 = (reg237 > reg224);
              reg254 <= ($unsigned($signed(((~|reg192) <= $signed(wire179)))) || ($signed(reg205) ?
                  (+reg207) : (|(~|(|(8'ha2))))));
            end
          else
            begin
              reg254 <= $unsigned($unsigned(($signed($unsigned(reg244)) >>> (reg236[(5'h15):(5'h10)] ?
                  (wire200 ? forvar239 : (8'hab)) : "R3"))));
              reg255 <= reg181;
            end
        end
      else
        begin
          reg247 = wire174;
          if ({(reg247 ?
                  $unsigned({(reg197 >> reg246)}) : (($unsigned(forvar232) ?
                          reg241[(4'hd):(3'h4)] : (reg204 ? wire177 : reg237)) ?
                      reg244 : forvar239[(3'h4):(1'h0)])),
              $signed($signed(reg204[(3'h5):(3'h4)]))})
            begin
              reg251 = (~^(~|wire179[(1'h1):(1'h1)]));
              reg254 <= reg248;
              reg255 <= $signed(reg183[(4'hb):(4'h8)]);
              reg256 <= reg191[(3'h4):(3'h4)];
              reg257 <= ($signed((reg218[(1'h1):(1'h0)] ?
                      "FLzfcXPm2" : (8'h9f))) ?
                  $signed(reg241) : reg218[(4'ha):(4'h9)]);
            end
          else
            begin
              reg248 <= {((~reg198[(4'h9):(3'h4)]) < {"AFBd1Mk4nxVz"})};
              reg249 <= reg197[(3'h4):(1'h1)];
              reg250 <= (|"TJeW4BToIkMGobt");
              reg251 = ($unsigned(((!(8'ha6)) <= reg242[(1'h1):(1'h0)])) ^ reg240[(3'h4):(1'h1)]);
              reg254 <= (reg205 != reg255[(3'h5):(2'h3)]);
            end
          for (forvar258 = (1'h0); (forvar258 < (1'h0)); forvar258 = (forvar258 + (1'h1)))
            begin
              reg259 = (!$signed(($signed((|reg238)) | reg209)));
              reg260 <= (&$signed(((wire173 <<< {reg230}) ?
                  (~(!reg182)) : $signed(wire174[(2'h2):(2'h2)]))));
              reg261 <= ("GQvomPvbk4sseKKy" ?
                  (wire200[(3'h6):(1'h0)] ?
                      $signed(reg230[(1'h0):(1'h0)]) : $signed((wire177 ?
                          (reg249 ?
                              reg181 : reg205) : $signed(reg256)))) : (8'hab));
              reg262 <= "";
              reg263 = ({((|$unsigned(reg214)) ?
                      $signed((reg229 ?
                          reg218 : wire177)) : (~|$signed(reg197))),
                  reg197[(2'h2):(1'h0)]} < (+((+$unsigned(reg198)) ?
                  ((~|reg233) ?
                      $unsigned(reg262) : $signed(reg260)) : $signed("JtyrnosyUp"))));
            end
          if ($unsigned((+$signed(((~(8'hb2)) * reg244[(3'h6):(1'h0)])))))
            begin
              reg264 <= (reg237[(2'h3):(2'h2)] & $signed(reg219[(1'h0):(1'h0)]));
              reg265 <= (reg257[(5'h12):(4'hf)] <<< $signed({(&$signed(reg238)),
                  $unsigned((wire174 * reg224))}));
              reg266 <= (reg259 ?
                  $unsigned($unsigned($unsigned($unsigned(reg183)))) : forvar232);
              reg267 <= reg209;
              reg268 <= $signed($signed(reg209[(4'hc):(4'ha)]));
            end
          else
            begin
              reg264 <= reg244[(3'h7):(2'h2)];
              reg265 <= reg230[(1'h0):(1'h0)];
              reg266 <= (!reg240);
            end
        end
      reg269 = $unsigned(reg235);
    end
  always
    @(posedge clk) begin
      reg270 <= ((|((8'ha3) + {(~reg246),
          (reg192 ? reg207 : wire174)})) == reg183);
      reg271 <= (reg262[(1'h1):(1'h0)] ?
          (reg243 <= (&(reg233[(5'h12):(5'h12)] ?
              $signed(wire199) : {reg219}))) : (|($signed(wire200) ?
              wire201 : (^~reg254[(1'h1):(1'h0)]))));
      reg272 <= $signed($unsigned(reg198[(1'h1):(1'h0)]));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module65
#(parameter param165 = {((+(8'hab)) ? (8'hbb) : {(^(^~(7'h44))), {((8'hb1) ? (8'hbe) : (8'hb7)), {(8'ha6), (8'hab)}}}), (^~{((^~(8'ha9)) > {(8'ha1)}), {(8'hb5), ((8'hb8) << (8'h9e))}})}, 
parameter param166 = (-{(8'hbb), (+param165)}))
(y, clk, wire70, wire69, wire68, wire67, wire66);
  output wire [(32'h474):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire70;
  input wire signed [(3'h7):(1'h0)] wire69;
  input wire signed [(4'hf):(1'h0)] wire68;
  input wire signed [(4'h9):(1'h0)] wire67;
  input wire [(5'h13):(1'h0)] wire66;
  wire signed [(5'h14):(1'h0)] wire164;
  wire [(4'ha):(1'h0)] wire150;
  wire signed [(4'hf):(1'h0)] wire119;
  wire signed [(5'h14):(1'h0)] wire118;
  wire [(4'hd):(1'h0)] wire117;
  wire [(5'h13):(1'h0)] wire116;
  wire signed [(4'hd):(1'h0)] wire115;
  wire signed [(4'hd):(1'h0)] wire114;
  wire signed [(3'h7):(1'h0)] wire113;
  wire [(4'h9):(1'h0)] wire112;
  wire [(4'h9):(1'h0)] wire111;
  wire [(2'h2):(1'h0)] wire110;
  wire [(5'h14):(1'h0)] wire109;
  wire [(4'h9):(1'h0)] wire108;
  wire signed [(5'h10):(1'h0)] wire107;
  wire [(2'h3):(1'h0)] wire105;
  wire [(5'h13):(1'h0)] wire84;
  reg [(4'hd):(1'h0)] reg161 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg160 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg159 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg156 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg155 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg152 = (1'h0);
  reg [(5'h12):(1'h0)] reg147 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg146 = (1'h0);
  reg [(5'h14):(1'h0)] reg145 = (1'h0);
  reg [(4'hc):(1'h0)] reg143 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg139 = (1'h0);
  reg [(4'hf):(1'h0)] reg138 = (1'h0);
  reg [(5'h10):(1'h0)] reg137 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg132 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg131 = (1'h0);
  reg [(4'ha):(1'h0)] reg130 = (1'h0);
  reg [(4'hc):(1'h0)] reg128 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg127 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg126 = (1'h0);
  reg [(4'hf):(1'h0)] reg123 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg122 = (1'h0);
  reg [(3'h5):(1'h0)] reg106 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg100 = (1'h0);
  reg [(4'h8):(1'h0)] reg98 = (1'h0);
  reg [(4'hc):(1'h0)] reg97 = (1'h0);
  reg [(4'hf):(1'h0)] reg94 = (1'h0);
  reg [(2'h2):(1'h0)] reg93 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg89 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg87 = (1'h0);
  reg [(4'h8):(1'h0)] reg83 = (1'h0);
  reg [(4'h8):(1'h0)] reg81 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg72 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg79 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg78 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg75 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg74 = (1'h0);
  reg [(5'h10):(1'h0)] reg71 = (1'h0);
  reg [(3'h5):(1'h0)] reg163 = (1'h0);
  reg [(2'h2):(1'h0)] reg162 = (1'h0);
  reg [(3'h5):(1'h0)] forvar158 = (1'h0);
  reg [(4'he):(1'h0)] reg157 = (1'h0);
  reg [(4'hd):(1'h0)] reg154 = (1'h0);
  reg [(5'h10):(1'h0)] reg153 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg151 = (1'h0);
  reg [(5'h14):(1'h0)] reg149 = (1'h0);
  reg [(5'h14):(1'h0)] reg148 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar144 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg142 = (1'h0);
  reg [(4'h9):(1'h0)] reg141 = (1'h0);
  reg [(5'h11):(1'h0)] forvar140 = (1'h0);
  reg [(5'h14):(1'h0)] reg136 = (1'h0);
  reg [(2'h3):(1'h0)] forvar135 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar134 = (1'h0);
  reg [(5'h10):(1'h0)] reg133 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar129 = (1'h0);
  reg [(5'h12):(1'h0)] reg125 = (1'h0);
  reg [(4'ha):(1'h0)] forvar124 = (1'h0);
  reg signed [(4'he):(1'h0)] reg121 = (1'h0);
  reg [(5'h12):(1'h0)] forvar120 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg104 = (1'h0);
  reg [(5'h13):(1'h0)] reg103 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar99 = (1'h0);
  reg [(5'h12):(1'h0)] forvar96 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg95 = (1'h0);
  reg [(5'h10):(1'h0)] reg92 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg91 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar90 = (1'h0);
  reg [(5'h10):(1'h0)] forvar88 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar86 = (1'h0);
  reg [(4'he):(1'h0)] reg85 = (1'h0);
  reg [(5'h13):(1'h0)] reg82 = (1'h0);
  reg [(2'h2):(1'h0)] reg80 = (1'h0);
  reg [(5'h12):(1'h0)] reg77 = (1'h0);
  reg [(5'h10):(1'h0)] forvar77 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg76 = (1'h0);
  reg [(2'h3):(1'h0)] reg73 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar72 = (1'h0);
  assign y = {wire164,
                 wire150,
                 wire119,
                 wire118,
                 wire117,
                 wire116,
                 wire115,
                 wire114,
                 wire113,
                 wire112,
                 wire111,
                 wire110,
                 wire109,
                 wire108,
                 wire107,
                 wire105,
                 wire84,
                 reg161,
                 reg160,
                 reg159,
                 reg156,
                 reg155,
                 reg152,
                 reg147,
                 reg146,
                 reg145,
                 reg143,
                 reg139,
                 reg138,
                 reg137,
                 reg132,
                 reg131,
                 reg130,
                 reg128,
                 reg127,
                 reg126,
                 reg123,
                 reg122,
                 reg106,
                 reg102,
                 reg100,
                 reg98,
                 reg97,
                 reg94,
                 reg93,
                 reg89,
                 reg87,
                 reg83,
                 reg81,
                 reg72,
                 reg79,
                 reg78,
                 reg75,
                 reg74,
                 reg71,
                 reg163,
                 reg162,
                 forvar158,
                 reg157,
                 reg154,
                 reg153,
                 reg151,
                 reg149,
                 reg148,
                 forvar144,
                 reg142,
                 reg141,
                 forvar140,
                 reg136,
                 forvar135,
                 forvar134,
                 reg133,
                 forvar129,
                 reg125,
                 forvar124,
                 reg121,
                 forvar120,
                 reg104,
                 reg103,
                 reg101,
                 forvar99,
                 forvar96,
                 reg95,
                 reg92,
                 reg91,
                 forvar90,
                 forvar88,
                 forvar86,
                 reg85,
                 reg82,
                 reg80,
                 reg77,
                 forvar77,
                 reg76,
                 reg73,
                 forvar72,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg71 <= (^(~&(|wire69)));
      if (reg71)
        begin
          for (forvar72 = (1'h0); (forvar72 < (3'h4)); forvar72 = (forvar72 + (1'h1)))
            begin
              reg73 = ("tTnTRT" <= wire66[(4'hc):(3'h7)]);
              reg74 <= reg71;
            end
          reg75 <= (~|$signed((&({wire66, (8'hbf)} ?
              (reg71 || (8'hbd)) : $unsigned(reg71)))));
          reg76 = ((~|(~&forvar72[(1'h0):(1'h0)])) + (~&$signed($unsigned((&reg71)))));
          for (forvar77 = (1'h0); (forvar77 < (1'h0)); forvar77 = (forvar77 + (1'h1)))
            begin
              reg78 <= {$unsigned((reg76 ?
                      (wire69[(1'h0):(1'h0)] ^ $signed((8'hac))) : (~|{reg71}))),
                  ($unsigned($unsigned(reg75[(2'h2):(2'h2)])) >= (reg74[(2'h3):(2'h2)] ?
                      ((wire70 ? forvar72 : reg74) ?
                          (wire66 ?
                              (8'hb8) : wire68) : (reg75 & reg76)) : reg74))};
              reg79 <= reg76;
            end
        end
      else
        begin
          if ({$signed(({$signed((8'had)), "P0GoSxvoE"} ?
                  reg78[(4'hf):(2'h2)] : $unsigned($unsigned(forvar77))))})
            begin
              reg72 <= wire70;
              reg73 = (wire67 ?
                  $unsigned(wire66[(4'hd):(4'ha)]) : $signed((7'h44)));
              reg76 = wire66;
              reg77 = reg72[(2'h3):(2'h3)];
              reg78 <= (wire69[(1'h0):(1'h0)] > $signed({({forvar77,
                      wire67} != $unsigned(wire70)),
                  $signed($unsigned(reg77))}));
            end
          else
            begin
              reg72 <= (reg76 != (+{$unsigned((forvar72 < reg78))}));
              reg74 <= ((-((reg77 ^ $signed(reg77)) <<< $signed("LWg7yMRG60SFBg9S"))) ?
                  $unsigned(reg78[(3'h5):(3'h4)]) : ($unsigned($signed(wire66)) | (~($signed(forvar77) ?
                      (reg76 ? reg76 : wire67) : (reg71 ~^ reg72)))));
            end
          reg80 = $signed(wire66[(1'h1):(1'h0)]);
        end
      reg81 <= reg79[(3'h4):(2'h3)];
      reg82 = wire69;
      reg83 <= (reg76[(2'h3):(1'h1)] ?
          {{((reg73 >= (8'hb5)) ? $unsigned(forvar72) : (8'hbe))},
              $unsigned(((!wire68) ?
                  "iHMZ3iKDM" : $signed(wire66)))} : ((($unsigned(forvar72) ?
              ((8'ha8) ?
                  reg82 : (7'h42)) : (|wire67)) >> wire67) + {($signed(reg72) >= (+wire67)),
              reg82[(4'hc):(4'h8)]}));
    end
  assign wire84 = {reg83, wire69};
  always
    @(posedge clk) begin
      reg85 = $signed(reg72);
      for (forvar86 = (1'h0); (forvar86 < (2'h2)); forvar86 = (forvar86 + (1'h1)))
        begin
          reg87 <= reg79[(1'h0):(1'h0)];
        end
      for (forvar88 = (1'h0); (forvar88 < (1'h0)); forvar88 = (forvar88 + (1'h1)))
        begin
          reg89 <= ({(reg79[(3'h7):(2'h3)] ?
                  (8'ha2) : $signed((wire68 ? wire69 : reg87))),
              $unsigned((reg74[(3'h4):(3'h4)] >>> $unsigned(forvar86)))} | (&(|{wire69})));
          for (forvar90 = (1'h0); (forvar90 < (1'h1)); forvar90 = (forvar90 + (1'h1)))
            begin
              reg91 = (-wire68[(4'ha):(3'h7)]);
              reg92 = (reg89[(3'h4):(1'h0)] || $signed(wire66));
              reg93 <= reg79;
              reg94 <= (reg79 ?
                  ($signed("rdvkKWNetOkJ") ?
                      reg87 : ((&reg89) <= (forvar88[(5'h10):(3'h5)] ?
                          $signed(reg79) : (reg93 ?
                              (8'haf) : reg74)))) : wire84);
              reg95 = reg91[(4'h9):(2'h2)];
            end
        end
      for (forvar96 = (1'h0); (forvar96 < (2'h3)); forvar96 = (forvar96 + (1'h1)))
        begin
          reg97 <= {$signed((~^({wire69} >= reg83[(3'h7):(3'h5)])))};
          reg98 <= ($signed((8'haf)) ?
              (~|$unsigned($unsigned(forvar96))) : (^(~|("n" ?
                  (wire66 && (7'h41)) : ((7'h43) ? reg97 : forvar96)))));
          for (forvar99 = (1'h0); (forvar99 < (3'h4)); forvar99 = (forvar99 + (1'h1)))
            begin
              reg100 <= (8'hb2);
              reg101 = (+wire68[(3'h4):(1'h0)]);
              reg102 <= reg83;
              reg103 = wire67[(1'h0):(1'h0)];
              reg104 = {$unsigned((~|($signed((8'h9f)) ?
                      (|reg75) : (|reg91))))};
            end
        end
    end
  assign wire105 = ({{wire84[(1'h0):(1'h0)]}, "7i"} ?
                       $unsigned(reg72[(1'h1):(1'h0)]) : $unsigned($signed({(+reg71),
                           $unsigned((8'hba))})));
  always
    @(posedge clk) begin
      reg106 <= $signed(reg93);
    end
  assign wire107 = $unsigned(reg97[(3'h5):(3'h4)]);
  assign wire108 = reg98[(1'h1):(1'h0)];
  assign wire109 = (8'ha3);
  assign wire110 = ($signed(((+(wire67 ?
                           wire108 : wire66)) || $signed(reg89))) ?
                       ($unsigned(reg81) ?
                           (($unsigned((8'hbb)) ?
                                   wire66 : (wire69 ? wire69 : reg94)) ?
                               $signed($unsigned(wire69)) : {$signed(reg97)}) : $unsigned({$unsigned(wire107)})) : $unsigned(((!(reg75 ?
                           (8'ha1) : reg97)) && $signed((^reg72)))));
  assign wire111 = (reg97 ?
                       reg79[(3'h4):(1'h1)] : $unsigned((~&"6p5KxVpKYKVeIfMfO5")));
  assign wire112 = ("h709QBr9VXSfED10zb" ?
                       "UR4hgiWAG7veSt2V6" : ($unsigned(((reg75 ^ reg100) ?
                           $signed(wire69) : $signed(reg83))) < $signed(((reg89 ^~ wire109) != ((8'hb4) >= reg71)))));
  assign wire113 = $signed(reg81[(3'h4):(1'h1)]);
  assign wire114 = ($signed((&((wire69 ? (8'ha8) : wire110) >= (~|reg78)))) ?
                       (reg71 <= (^~(reg74[(4'ha):(2'h3)] ?
                           $signed((8'h9c)) : $signed(reg102)))) : wire112[(3'h4):(1'h0)]);
  assign wire115 = (8'h9c);
  assign wire116 = {$unsigned((($unsigned(reg72) ? $signed(reg72) : (|wire67)) ?
                           $unsigned((wire115 != wire107)) : ({(7'h43),
                               reg87} || $unsigned(reg106))))};
  assign wire117 = $signed($unsigned(((&(wire110 ?
                       reg98 : reg93)) && $signed((~(7'h43))))));
  assign wire118 = {{(^~wire70[(3'h4):(2'h3)])}, "YqlVd8xO1YI3wPL1hJBV"};
  assign wire119 = ((-{((reg87 >>> reg87) <= $unsigned(wire107))}) - $signed(reg79));
  always
    @(posedge clk) begin
      for (forvar120 = (1'h0); (forvar120 < (1'h0)); forvar120 = (forvar120 + (1'h1)))
        begin
          reg121 = (((~$signed(reg100)) >= reg98) ?
              reg87[(1'h1):(1'h1)] : (!($signed($unsigned(wire118)) >= $unsigned(reg83[(1'h0):(1'h0)]))));
          reg122 <= ($unsigned($signed((&wire111[(2'h3):(1'h1)]))) ?
              (^~$unsigned((((7'h44) ? reg81 : (8'hbc)) ?
                  (&reg89) : $unsigned(wire116)))) : (($unsigned($unsigned(reg81)) ?
                      $signed("Hyl7RI9Ons") : $signed((|wire108))) ?
                  (((wire84 ?
                      wire110 : wire68) >>> $unsigned(wire116)) >> reg83) : reg87));
          reg123 <= (~&"HDbhPAArQgVd1Y");
          for (forvar124 = (1'h0); (forvar124 < (1'h1)); forvar124 = (forvar124 + (1'h1)))
            begin
              reg125 = (~&(8'ha2));
              reg126 <= {wire117[(4'hb):(1'h0)],
                  {"qZDf9WWEGLes5s", {wire67, (~|(reg93 && reg87))}}};
              reg127 <= (((reg74[(3'h6):(3'h4)] << ("Js2oxs9" ?
                      $signed(reg123) : $unsigned(reg122))) == "x4b13zHcbr") ?
                  (~&(reg123 && $signed((&reg81)))) : $unsigned(($unsigned($unsigned(reg123)) + reg97)));
              reg128 <= ({$signed((((8'hb3) ? wire70 : wire113) ?
                      $signed(wire114) : reg123))} == $unsigned((~&$signed(((8'hb0) >> wire69)))));
            end
          for (forvar129 = (1'h0); (forvar129 < (2'h3)); forvar129 = (forvar129 + (1'h1)))
            begin
              reg130 <= "h9LNkYvioddSPxiODFEz";
              reg131 <= wire66;
              reg132 <= (8'ha1);
            end
        end
      reg133 = (~|(|$unsigned((^~reg87[(2'h2):(2'h2)]))));
      for (forvar134 = (1'h0); (forvar134 < (1'h1)); forvar134 = (forvar134 + (1'h1)))
        begin
          for (forvar135 = (1'h0); (forvar135 < (1'h1)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 = ($signed({(&$unsigned(reg131)), reg72}) ?
                  forvar134 : {(forvar129 ?
                          {reg71[(1'h1):(1'h1)]} : ($signed((8'ha4)) == (reg123 ?
                              (8'ha4) : reg126)))});
              reg137 <= (|($unsigned(wire68[(3'h5):(1'h0)]) == $signed({(reg100 - reg127),
                  wire108})));
              reg138 <= $signed({($signed((reg83 >= wire69)) & {(wire114 ?
                          wire108 : (8'hac))}),
                  {($unsigned(wire111) ?
                          "qbfaimNLe4Bag9qrihCZ" : (wire118 ~^ forvar120))}});
              reg139 <= ((($signed($signed(reg72)) ?
                          reg98 : $unsigned($signed(reg122))) ?
                      $signed((forvar124 != (wire118 ?
                          reg75 : reg126))) : ($unsigned((reg98 ?
                          reg123 : wire66)) ^ {(-(8'hbc))})) ?
                  $unsigned((reg89 || $signed((wire112 - reg126)))) : (-$signed(((^reg132) <<< reg102))));
            end
          for (forvar140 = (1'h0); (forvar140 < (3'h4)); forvar140 = (forvar140 + (1'h1)))
            begin
              reg141 = (^~(reg98 ? $signed((^reg123)) : reg132));
              reg142 = (~^(reg123 ?
                  {reg133[(2'h3):(2'h2)],
                      (reg106 == (~|reg131))} : ($unsigned($unsigned(wire109)) + wire119)));
            end
          reg143 <= wire67[(4'h8):(1'h1)];
        end
      for (forvar144 = (1'h0); (forvar144 < (3'h4)); forvar144 = (forvar144 + (1'h1)))
        begin
          if ((&forvar124[(2'h3):(1'h1)]))
            begin
              reg145 <= wire110;
              reg146 <= wire105;
              reg147 <= $unsigned((forvar129[(3'h7):(2'h3)] ?
                  {((reg146 >>> reg143) ?
                          {wire69} : "WtnY6ewRGTL6ro")} : $unsigned(({reg93} ?
                      (reg133 ? (8'hb0) : reg128) : $unsigned(wire117)))));
            end
          else
            begin
              reg148 = (^(reg139 ?
                  "q9is5TzEX7" : ($unsigned($unsigned(wire113)) ?
                      ($unsigned(wire117) | (+forvar129)) : "lOHL70LeYv5Mqsw")));
              reg149 = $signed((({reg98[(1'h0):(1'h0)]} ?
                      (^(reg145 ? reg126 : reg147)) : reg102) ?
                  $unsigned((!reg145[(5'h14):(3'h6)])) : $signed($unsigned($signed(reg127)))));
            end
        end
    end
  assign wire150 = $signed(($signed((7'h40)) << {$unsigned((reg106 ?
                           wire111 : reg146)),
                       $signed(wire118[(2'h3):(2'h3)])}));
  always
    @(posedge clk) begin
      if ((^~(^~$signed(reg102[(2'h3):(2'h2)]))))
        begin
          if (($unsigned("BEX3M6HWOttw") ?
              $unsigned($unsigned(reg123)) : $signed({reg89[(1'h1):(1'h1)]})))
            begin
              reg151 = $unsigned($signed(($unsigned($signed(reg102)) ?
                  ({wire111} * wire116) : (wire117[(3'h6):(2'h2)] ?
                      reg83 : reg89))));
              reg152 <= (&reg71[(4'hc):(4'h9)]);
              reg153 = (~wire112);
              reg154 = (&(wire107[(3'h5):(2'h3)] ^ (reg128 + $unsigned($signed(reg93)))));
              reg155 <= $unsigned(wire70);
            end
          else
            begin
              reg151 = (8'ha8);
              reg152 <= (^~wire117);
            end
        end
      else
        begin
          reg152 <= $unsigned($signed($unsigned(($signed(wire113) && $unsigned(wire68)))));
          if ((^wire119))
            begin
              reg155 <= $signed((|{$signed((wire67 ? (8'ha4) : reg93))}));
              reg156 <= (+"uE");
            end
          else
            begin
              reg155 <= {"cyCLd46hCuo49YlllHi"};
              reg157 = (wire110 ? wire105[(2'h3):(1'h1)] : wire114);
            end
          for (forvar158 = (1'h0); (forvar158 < (3'h4)); forvar158 = (forvar158 + (1'h1)))
            begin
              reg159 <= $unsigned($unsigned($signed(((reg152 ?
                      wire66 : reg157) ?
                  (reg154 ? (8'hb4) : reg72) : $signed(reg130)))));
              reg160 <= {reg79};
              reg161 <= $signed(reg153[(4'hb):(2'h3)]);
              reg162 = {$unsigned((|$signed((reg131 ? reg130 : reg159)))),
                  {$unsigned((reg143[(2'h3):(2'h3)] ^~ {(8'haa)})),
                      wire115[(2'h3):(1'h1)]}};
            end
          reg163 = (wire150[(2'h2):(1'h0)] | reg87[(1'h0):(1'h0)]);
        end
    end
  assign wire164 = (reg123[(4'hf):(4'he)] ?
                       reg74 : $unsigned(reg97[(4'hc):(3'h4)]));
endmodule