(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h84):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire0;
  input wire [(5'h14):(1'h0)] wire1;
  input wire [(4'he):(1'h0)] wire2;
  input wire signed [(5'h12):(1'h0)] wire3;
  wire signed [(2'h3):(1'h0)] wire442;
  wire [(4'hc):(1'h0)] wire440;
  wire signed [(4'he):(1'h0)] wire439;
  wire [(2'h2):(1'h0)] wire438;
  wire [(4'hb):(1'h0)] wire437;
  wire signed [(4'he):(1'h0)] wire436;
  wire signed [(4'h9):(1'h0)] wire435;
  wire [(4'hc):(1'h0)] wire4;
  wire signed [(5'h15):(1'h0)] wire5;
  wire [(5'h15):(1'h0)] wire6;
  wire signed [(4'hc):(1'h0)] wire433;
  assign y = {wire442,
                 wire440,
                 wire439,
                 wire438,
                 wire437,
                 wire436,
                 wire435,
                 wire4,
                 wire5,
                 wire6,
                 wire433,
                 (1'h0)};
  assign wire4 = wire1;
  assign wire5 = (wire1 <= ($signed(((wire3 ? wire1 : wire3) ^ ((8'ha3) ?
                         wire4 : wire0))) ?
                     wire2[(1'h1):(1'h0)] : $unsigned(wire4)));
  assign wire6 = wire1;
  module7 #() modinst434 (.wire11(wire1), .clk(clk), .wire12(wire0), .wire8(wire4), .wire9(wire5), .wire10(wire6), .y(wire433));
  assign wire435 = ({wire5, wire6} - wire433);
  assign wire436 = ((~^wire435[(3'h6):(3'h4)]) ?
                       wire6 : ((~&(wire3 ?
                           (wire0 ^ wire3) : {wire433})) ~^ $signed(($signed((7'h41)) | wire2[(1'h0):(1'h0)]))));
  assign wire437 = wire3;
  assign wire438 = $signed($unsigned((({wire6, wire2} ?
                           wire4[(4'ha):(3'h5)] : $unsigned((8'h9e))) ?
                       wire2 : ((+wire435) | (wire6 >> wire4)))));
  assign wire439 = (+(({(8'hbe), $unsigned((8'ha0))} ?
                       (~|$signed(wire436)) : (wire438 ?
                           $signed(wire2) : (wire437 ^ wire5))) == (wire436[(2'h2):(1'h0)] ?
                       {$signed(wire6)} : (wire5[(5'h15):(5'h11)] >= wire3[(3'h4):(3'h4)]))));

  assign wire442 = $unsigned((!(((wire5 ?
                       wire2 : wire437) >= (~^wire435)) >>> ($signed(wire0) == (wire2 > wire2)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module7  (y, clk, wire12, wire11, wire10, wire9, wire8);
  output wire [(32'hc6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire12;
  input wire [(5'h14):(1'h0)] wire11;
  input wire [(5'h15):(1'h0)] wire10;
  input wire signed [(5'h15):(1'h0)] wire9;
  input wire [(4'hc):(1'h0)] wire8;
  wire signed [(3'h6):(1'h0)] wire432;
  wire signed [(4'h9):(1'h0)] wire431;
  wire signed [(2'h2):(1'h0)] wire199;
  wire signed [(4'he):(1'h0)] wire91;
  wire signed [(5'h12):(1'h0)] wire89;
  wire signed [(4'he):(1'h0)] wire16;
  wire [(5'h14):(1'h0)] wire15;
  wire [(4'hd):(1'h0)] wire14;
  wire signed [(4'hb):(1'h0)] wire13;
  wire signed [(4'hc):(1'h0)] wire201;
  wire signed [(4'hb):(1'h0)] wire202;
  wire [(4'hc):(1'h0)] wire302;
  wire signed [(5'h12):(1'h0)] wire304;
  wire signed [(4'hf):(1'h0)] wire323;
  wire signed [(3'h4):(1'h0)] wire325;
  wire [(3'h7):(1'h0)] wire326;
  wire signed [(4'hb):(1'h0)] wire429;
  assign y = {wire432,
                 wire431,
                 wire199,
                 wire91,
                 wire89,
                 wire16,
                 wire15,
                 wire14,
                 wire13,
                 wire201,
                 wire202,
                 wire302,
                 wire304,
                 wire323,
                 wire325,
                 wire326,
                 wire429,
                 (1'h0)};
  assign wire13 = (^{$unsigned({(wire8 < wire8)})});
  assign wire14 = ((~(wire11[(1'h1):(1'h1)] ?
                      ($unsigned(wire12) ?
                          wire12[(4'hc):(4'ha)] : $signed(wire12)) : (!$signed(wire11)))) >> ($unsigned($signed((wire12 << (8'haf)))) != wire9));
  assign wire15 = $signed($signed($unsigned((((8'ha1) == wire14) & (7'h40)))));
  assign wire16 = ({(((~|wire9) ?
                              (wire13 ?
                                  wire11 : wire14) : wire11[(2'h3):(2'h2)]) & wire9)} ?
                      wire11[(3'h7):(3'h7)] : $signed({($signed(wire15) <<< (8'hb9)),
                          wire10[(4'hf):(3'h5)]}));

  assign wire91 = wire11;
  assign wire201 = (|wire9);
  assign wire202 = (&($unsigned($signed($signed(wire199))) ?
                       $unsigned($signed((wire91 ?
                           wire11 : wire91))) : (-wire13)));
  module203 #() modinst303 (.y(wire302), .wire205(wire202), .wire207(wire8), .clk(clk), .wire204(wire9), .wire206(wire13));
  assign wire304 = $unsigned(wire13[(3'h5):(3'h4)]);
  assign wire325 = (8'hbe);
  assign wire326 = (wire201[(3'h7):(3'h6)] ^ ((8'ha9) || (+(~(wire14 ^ wire8)))));
  assign wire431 = $unsigned(wire325);
  assign wire432 = $unsigned((+$signed($unsigned((wire431 ?
                       (8'hbf) : wire11)))));
endmodule



(* use_dsp48="no" *) (* use_dsp="no" *) module module203  (y, clk, wire207, wire206, wire205, wire204);
  output wire [(32'h45e):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire207;
  input wire [(4'h8):(1'h0)] wire206;
  input wire signed [(4'ha):(1'h0)] wire205;
  input wire [(5'h14):(1'h0)] wire204;
  wire signed [(4'hb):(1'h0)] wire301;
  wire [(4'hd):(1'h0)] wire300;
  wire signed [(4'hb):(1'h0)] wire299;
  wire [(5'h11):(1'h0)] wire298;
  wire [(5'h13):(1'h0)] wire297;
  wire [(5'h10):(1'h0)] wire296;
  wire signed [(3'h5):(1'h0)] wire295;
  wire signed [(5'h12):(1'h0)] wire294;
  wire [(4'h8):(1'h0)] wire293;
  wire signed [(4'hc):(1'h0)] wire292;
  wire signed [(4'ha):(1'h0)] wire291;
  wire [(4'h8):(1'h0)] wire277;
  wire signed [(5'h12):(1'h0)] wire276;
  wire signed [(3'h7):(1'h0)] wire275;
  wire [(5'h13):(1'h0)] wire274;
  wire [(5'h11):(1'h0)] wire273;
  reg signed [(4'ha):(1'h0)] reg290 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg288 = (1'h0);
  reg [(3'h6):(1'h0)] reg287 = (1'h0);
  reg [(4'ha):(1'h0)] reg286 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg285 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg283 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg282 = (1'h0);
  reg [(4'ha):(1'h0)] reg280 = (1'h0);
  reg signed [(4'he):(1'h0)] reg279 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg278 = (1'h0);
  reg [(4'hf):(1'h0)] reg272 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg271 = (1'h0);
  reg [(5'h15):(1'h0)] reg268 = (1'h0);
  reg [(5'h11):(1'h0)] reg267 = (1'h0);
  reg [(5'h10):(1'h0)] reg266 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg265 = (1'h0);
  reg [(3'h4):(1'h0)] reg262 = (1'h0);
  reg [(2'h2):(1'h0)] reg260 = (1'h0);
  reg [(3'h4):(1'h0)] reg256 = (1'h0);
  reg [(4'h8):(1'h0)] reg255 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg251 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg249 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg246 = (1'h0);
  reg [(4'hf):(1'h0)] reg243 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg240 = (1'h0);
  reg [(5'h11):(1'h0)] reg239 = (1'h0);
  reg [(3'h4):(1'h0)] reg236 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg235 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg231 = (1'h0);
  reg [(4'ha):(1'h0)] reg230 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg229 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg225 = (1'h0);
  reg [(5'h10):(1'h0)] reg224 = (1'h0);
  reg [(4'hd):(1'h0)] reg223 = (1'h0);
  reg [(4'ha):(1'h0)] reg222 = (1'h0);
  reg [(5'h13):(1'h0)] reg221 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg218 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg213 = (1'h0);
  reg [(4'hc):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar289 = (1'h0);
  reg [(5'h10):(1'h0)] forvar284 = (1'h0);
  reg [(2'h2):(1'h0)] reg281 = (1'h0);
  reg [(4'ha):(1'h0)] forvar278 = (1'h0);
  reg [(5'h13):(1'h0)] reg270 = (1'h0);
  reg [(5'h10):(1'h0)] forvar269 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar264 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg263 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg261 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg259 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar258 = (1'h0);
  reg [(3'h7):(1'h0)] reg257 = (1'h0);
  reg [(5'h10):(1'h0)] reg254 = (1'h0);
  reg [(5'h10):(1'h0)] forvar253 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar252 = (1'h0);
  reg [(2'h3):(1'h0)] reg250 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar248 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg247 = (1'h0);
  reg [(3'h6):(1'h0)] forvar245 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar244 = (1'h0);
  reg [(4'hd):(1'h0)] reg242 = (1'h0);
  reg [(5'h12):(1'h0)] reg241 = (1'h0);
  reg [(3'h6):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar237 = (1'h0);
  reg [(5'h14):(1'h0)] forvar234 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar233 = (1'h0);
  reg [(5'h10):(1'h0)] reg232 = (1'h0);
  reg [(5'h11):(1'h0)] forvar228 = (1'h0);
  reg [(4'hd):(1'h0)] reg227 = (1'h0);
  reg [(4'hd):(1'h0)] forvar226 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar220 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar219 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg217 = (1'h0);
  reg [(5'h14):(1'h0)] reg216 = (1'h0);
  reg [(5'h15):(1'h0)] reg215 = (1'h0);
  reg [(4'ha):(1'h0)] forvar214 = (1'h0);
  reg [(5'h11):(1'h0)] forvar212 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar209 = (1'h0);
  reg [(5'h12):(1'h0)] forvar208 = (1'h0);
  assign y = {wire301,
                 wire300,
                 wire299,
                 wire298,
                 wire297,
                 wire296,
                 wire295,
                 wire294,
                 wire293,
                 wire292,
                 wire291,
                 wire277,
                 wire276,
                 wire275,
                 wire274,
                 wire273,
                 reg290,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg283,
                 reg282,
                 reg280,
                 reg279,
                 reg278,
                 reg272,
                 reg271,
                 reg268,
                 reg267,
                 reg266,
                 reg265,
                 reg262,
                 reg260,
                 reg256,
                 reg255,
                 reg251,
                 reg249,
                 reg246,
                 reg243,
                 reg240,
                 reg239,
                 reg236,
                 reg235,
                 reg231,
                 reg230,
                 reg229,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg218,
                 reg213,
                 reg211,
                 forvar289,
                 forvar284,
                 reg281,
                 forvar278,
                 reg270,
                 forvar269,
                 forvar264,
                 reg263,
                 reg261,
                 reg259,
                 forvar258,
                 reg257,
                 reg254,
                 forvar253,
                 forvar252,
                 reg250,
                 forvar248,
                 reg247,
                 forvar245,
                 forvar244,
                 reg242,
                 reg241,
                 reg238,
                 forvar237,
                 forvar234,
                 forvar233,
                 reg232,
                 forvar228,
                 reg227,
                 forvar226,
                 forvar220,
                 forvar219,
                 reg217,
                 reg216,
                 reg215,
                 forvar214,
                 forvar212,
                 reg210,
                 forvar209,
                 forvar208,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar208 = (1'h0); (forvar208 < (2'h3)); forvar208 = (forvar208 + (1'h1)))
        begin
          for (forvar209 = (1'h0); (forvar209 < (1'h1)); forvar209 = (forvar209 + (1'h1)))
            begin
              reg210 = {(|wire205[(4'h9):(4'h8)])};
              reg211 <= (+((8'haf) ^ $unsigned($signed((-reg210)))));
            end
          for (forvar212 = (1'h0); (forvar212 < (1'h0)); forvar212 = (forvar212 + (1'h1)))
            begin
              reg213 <= forvar209[(4'h8):(2'h3)];
            end
          for (forvar214 = (1'h0); (forvar214 < (2'h3)); forvar214 = (forvar214 + (1'h1)))
            begin
              reg215 = (~^{forvar209[(3'h7):(2'h3)]});
              reg216 = ((&(((reg213 ?
                      wire204 : reg215) ^ ((8'hb7) ^~ (8'ha1))) ^ forvar212[(4'he):(4'he)])) ?
                  wire204 : (~^(!forvar214)));
            end
          reg217 = $unsigned(($unsigned($signed(reg216[(4'hd):(1'h1)])) ?
              (~&(!(forvar209 ?
                  reg210 : (8'hb8)))) : $unsigned((~$unsigned(wire207)))));
          reg218 <= ($unsigned({((reg211 ? wire207 : wire204) ?
                  (forvar212 | wire205) : $unsigned(forvar209)),
              $unsigned($unsigned(forvar208))}) <= reg211);
        end
      for (forvar219 = (1'h0); (forvar219 < (3'h4)); forvar219 = (forvar219 + (1'h1)))
        begin
          for (forvar220 = (1'h0); (forvar220 < (1'h1)); forvar220 = (forvar220 + (1'h1)))
            begin
              reg221 <= forvar214;
              reg222 <= $signed(($signed($unsigned((~forvar208))) ?
                  $unsigned(($unsigned(wire204) ?
                      ((8'hbc) ?
                          reg210 : reg213) : {(8'h9f)})) : {((wire207 & forvar212) == (^~forvar209)),
                      (wire206 * (wire205 != wire206))}));
              reg223 <= $signed($unsigned(forvar220[(4'h9):(3'h5)]));
              reg224 <= (reg217 ?
                  ((~^({wire206, (7'h43)} ?
                      reg216 : $signed((7'h40)))) > reg218[(2'h2):(1'h1)]) : (((!$unsigned(reg215)) ?
                      (|(reg216 ?
                          reg217 : (8'ha6))) : $unsigned($signed(forvar208))) && $signed($signed(reg211))));
              reg225 <= reg216;
            end
          for (forvar226 = (1'h0); (forvar226 < (2'h3)); forvar226 = (forvar226 + (1'h1)))
            begin
              reg227 = reg224[(4'hd):(4'hb)];
            end
          for (forvar228 = (1'h0); (forvar228 < (1'h0)); forvar228 = (forvar228 + (1'h1)))
            begin
              reg229 <= forvar219;
              reg230 <= reg217[(3'h4):(2'h3)];
              reg231 <= {{forvar228[(4'h9):(2'h3)],
                      $unsigned(((|reg211) - $unsigned(reg217)))}};
            end
        end
      reg232 = $signed(reg229);
    end
  always
    @(posedge clk) begin
      for (forvar233 = (1'h0); (forvar233 < (2'h2)); forvar233 = (forvar233 + (1'h1)))
        begin
          for (forvar234 = (1'h0); (forvar234 < (2'h3)); forvar234 = (forvar234 + (1'h1)))
            begin
              reg235 <= wire204[(4'hd):(1'h0)];
              reg236 <= wire204[(1'h1):(1'h0)];
            end
          for (forvar237 = (1'h0); (forvar237 < (1'h1)); forvar237 = (forvar237 + (1'h1)))
            begin
              reg238 = ((reg224[(4'hd):(2'h3)] ?
                  (((^~reg218) ?
                      wire207 : (forvar233 ?
                          (7'h41) : reg213)) << $unsigned({reg211})) : ((+reg218) ?
                      (^~reg230[(4'ha):(3'h5)]) : $unsigned((forvar233 >> reg235)))) >> {(reg229[(2'h3):(2'h3)] ?
                      $signed((~^reg231)) : (~$signed(reg213)))});
              reg239 <= (~{(~&wire204[(5'h12):(3'h5)]), reg218});
              reg240 <= reg236[(3'h4):(1'h1)];
              reg241 = reg240;
              reg242 = (reg221 & wire204);
            end
          reg243 <= (($signed((8'ha4)) ?
                  (reg225 ?
                      reg230[(3'h4):(1'h1)] : $signed((reg236 <= wire205))) : $signed(wire204)) ?
              {(&(wire206 > {reg235}))} : (~{(|(reg213 ? reg240 : reg240)),
                  (&(reg230 ? wire207 : reg224))}));
        end
      for (forvar244 = (1'h0); (forvar244 < (3'h4)); forvar244 = (forvar244 + (1'h1)))
        begin
          for (forvar245 = (1'h0); (forvar245 < (1'h1)); forvar245 = (forvar245 + (1'h1)))
            begin
              reg246 <= ($unsigned(({$unsigned(forvar237),
                  $signed((8'ha8))} << {(-forvar244),
                  reg229})) <= $signed(reg241));
              reg247 = $unsigned($unsigned(($unsigned((reg243 >= wire206)) == (((7'h41) ?
                      reg243 : forvar237) ?
                  $unsigned(reg246) : (~&reg224)))));
            end
          for (forvar248 = (1'h0); (forvar248 < (2'h3)); forvar248 = (forvar248 + (1'h1)))
            begin
              reg249 <= (+reg240[(2'h2):(1'h1)]);
              reg250 = reg240[(4'h8):(2'h2)];
              reg251 <= ((forvar244[(2'h2):(1'h0)] ?
                      ($unsigned((~|reg242)) != (8'hbf)) : reg241) ?
                  ($unsigned((~&(reg223 ? reg247 : wire207))) ?
                      $signed((reg225 ?
                          {(8'hb9)} : $unsigned(reg235))) : wire205) : (reg211[(4'hc):(2'h2)] & reg231));
            end
        end
      for (forvar252 = (1'h0); (forvar252 < (1'h1)); forvar252 = (forvar252 + (1'h1)))
        begin
          for (forvar253 = (1'h0); (forvar253 < (2'h2)); forvar253 = (forvar253 + (1'h1)))
            begin
              reg254 = ($unsigned($unsigned($signed((7'h40)))) >> (8'ha0));
              reg255 <= reg222;
              reg256 <= $unsigned($unsigned({$unsigned((reg235 ?
                      reg211 : (8'hb4))),
                  reg243}));
              reg257 = reg218[(2'h3):(2'h2)];
            end
          for (forvar258 = (1'h0); (forvar258 < (2'h3)); forvar258 = (forvar258 + (1'h1)))
            begin
              reg259 = ((reg246 >>> (~&$unsigned({forvar234}))) || {$signed($unsigned((+forvar245)))});
              reg260 <= reg239;
              reg261 = reg222;
              reg262 <= (8'hbc);
              reg263 = (^~(~^(8'h9d)));
            end
          for (forvar264 = (1'h0); (forvar264 < (2'h3)); forvar264 = (forvar264 + (1'h1)))
            begin
              reg265 <= reg229[(2'h3):(2'h3)];
              reg266 <= $signed(forvar264[(1'h1):(1'h1)]);
              reg267 <= $signed($unsigned($unsigned($signed(wire206))));
              reg268 <= reg266[(3'h7):(2'h3)];
            end
          for (forvar269 = (1'h0); (forvar269 < (1'h1)); forvar269 = (forvar269 + (1'h1)))
            begin
              reg270 = $unsigned({$signed($signed($signed(reg223)))});
              reg271 <= $signed({{(|$unsigned(reg254))},
                  $unsigned({forvar253[(2'h3):(1'h0)],
                      reg240[(4'ha):(3'h7)]})});
              reg272 <= ($signed((^~($signed(reg257) ~^ (reg231 > forvar264)))) - ($signed($signed((~|reg257))) ?
                  (~|$unsigned($signed(wire206))) : reg265));
            end
        end
    end
  assign wire273 = (($signed($signed((~&reg223))) ?
                           {(&$unsigned((8'hb5))),
                               ((reg236 ? (8'ha0) : reg249) ?
                                   $signed(reg251) : reg243[(4'hf):(3'h4)])} : ({(!reg255),
                               $signed(reg266)} ~^ reg271)) ?
                       ({(reg222 | ((8'haa) ? (8'ha0) : reg246)),
                               (~$unsigned((8'ha2)))} ?
                           (^(~&(8'ha1))) : {reg239,
                               (&(8'ha5))}) : (reg267[(3'h7):(2'h3)] ?
                           $signed($signed((reg260 > reg222))) : $unsigned((~^(reg221 - reg267)))));
  assign wire274 = (wire273[(4'ha):(3'h5)] ?
                       (~|((reg271 ? reg222[(3'h6):(3'h5)] : wire207) ?
                           wire207 : (-$unsigned(reg268)))) : (8'ha6));
  assign wire275 = ((&$signed(reg249)) ? reg218[(2'h3):(1'h1)] : reg230);
  assign wire276 = reg229[(4'hd):(4'hd)];
  assign wire277 = $unsigned($signed(($unsigned((^wire275)) & ($signed((8'hb1)) ?
                       $signed(reg266) : {reg260, (8'hb8)}))));
  always
    @(posedge clk) begin
      if ((((~|$signed({reg218})) ^ ((+$signed(reg231)) ?
          reg255[(3'h6):(2'h3)] : (~|{(8'hb9)}))) | reg272[(4'h8):(3'h6)]))
        begin
          reg278 <= (^{$signed(reg236)});
          reg279 <= $signed(reg268);
        end
      else
        begin
          for (forvar278 = (1'h0); (forvar278 < (3'h4)); forvar278 = (forvar278 + (1'h1)))
            begin
              reg279 <= (($unsigned($signed($signed(reg260))) ?
                      $unsigned((+(-reg272))) : ($signed((~reg225)) - (reg222 <<< $signed((8'h9f))))) ?
                  ($unsigned({reg271[(3'h6):(1'h1)]}) - (~(reg262[(1'h0):(1'h0)] ?
                      (reg230 != reg279) : {wire207, wire275}))) : (8'ha9));
              reg280 <= reg236;
              reg281 = {(&reg260),
                  (-($signed((|reg223)) ?
                      {$signed(reg262)} : ((^(8'ha1)) ?
                          (wire277 ? reg246 : (8'hb1)) : $unsigned(reg266))))};
              reg282 <= $signed($unsigned($signed({(reg280 ?
                      reg249 : wire205)})));
            end
          reg283 <= {((8'ha7) ?
                  (~|((8'hb0) ? reg224 : (!wire277))) : {(8'ha5)}),
              ((^(+(^reg213))) ?
                  reg230[(3'h6):(3'h6)] : {reg239[(3'h6):(1'h0)]})};
          for (forvar284 = (1'h0); (forvar284 < (2'h2)); forvar284 = (forvar284 + (1'h1)))
            begin
              reg285 <= (~|wire273);
              reg286 <= reg283[(1'h0):(1'h0)];
              reg287 <= reg278;
              reg288 <= reg224;
            end
          for (forvar289 = (1'h0); (forvar289 < (1'h0)); forvar289 = (forvar289 + (1'h1)))
            begin
              reg290 <= ($unsigned({(~(^~reg213)),
                      $unsigned($unsigned(reg211))}) ?
                  $signed(({(~wire274), (reg282 != reg249)} ?
                      $signed((reg281 ?
                          reg225 : reg278)) : $unsigned(wire273))) : wire205);
            end
        end
    end
  assign wire291 = $signed($unsigned((|reg279)));
  assign wire292 = $signed((&(((wire205 || (8'hae)) ?
                           $unsigned((8'ha3)) : (+reg256)) ?
                       $signed($signed(reg246)) : (reg221[(4'hf):(4'hb)] ?
                           $unsigned(reg283) : (reg230 ? reg287 : reg256)))));
  assign wire293 = {$unsigned(reg287),
                       $signed($signed(((reg268 ? reg223 : reg290) ?
                           $unsigned(reg268) : {wire206, wire274})))};
  assign wire294 = (~reg230[(3'h7):(2'h3)]);
  assign wire295 = $unsigned(($signed(($signed(reg225) << (8'ha4))) + (~&(!$unsigned(wire206)))));
  assign wire296 = {$signed($unsigned((~$unsigned(reg265))))};
  assign wire297 = (reg255 <<< wire276[(4'he):(2'h2)]);
  assign wire298 = reg287[(1'h1):(1'h0)];
  assign wire299 = (wire205[(2'h3):(2'h2)] && {(~&reg246)});
  assign wire300 = (reg231[(2'h2):(2'h2)] > (wire275[(1'h1):(1'h0)] < wire204));
  assign wire301 = (^(reg211[(4'ha):(4'h9)] ?
                       (((reg290 ? (8'haf) : (8'hb0)) ^ wire292) ?
                           {wire204} : ($signed(reg229) ?
                               reg266[(1'h0):(1'h0)] : reg290)) : $signed($unsigned((~|reg239)))));
endmodule


