module top
#(parameter param226 = ({((&(7'h42)) && (8'hb5)), {({(8'had), (8'ha6)} ? (8'ha1) : ((7'h41) | (8'ha7)))}} ? (&(~&(((8'h9c) + (8'hb0)) ? ((8'haa) ? (8'h9c) : (8'hb7)) : (8'haa)))) : (8'hb7)), 
parameter param227 = {param226})
(y, clk, wire0, wire1, wire2, wire3, wire4);
  output wire [(32'h1e6):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h13):(1'h0)] wire0;
  input wire signed [(4'hd):(1'h0)] wire1;
  input wire [(5'h12):(1'h0)] wire2;
  input wire signed [(4'hb):(1'h0)] wire3;
  input wire signed [(4'h8):(1'h0)] wire4;
  wire [(5'h14):(1'h0)] wire225;
  wire signed [(2'h3):(1'h0)] wire224;
  wire signed [(4'ha):(1'h0)] wire187;
  reg [(4'hc):(1'h0)] reg223 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg220 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg219 = (1'h0);
  reg [(5'h12):(1'h0)] reg217 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg216 = (1'h0);
  reg [(4'h9):(1'h0)] reg215 = (1'h0);
  reg [(4'h9):(1'h0)] reg211 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg209 = (1'h0);
  reg [(5'h15):(1'h0)] reg208 = (1'h0);
  reg [(2'h2):(1'h0)] reg207 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg206 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg205 = (1'h0);
  reg [(2'h3):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg203 = (1'h0);
  reg [(5'h15):(1'h0)] reg202 = (1'h0);
  reg [(5'h11):(1'h0)] reg201 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg199 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg198 = (1'h0);
  reg [(3'h7):(1'h0)] reg197 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg196 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg195 = (1'h0);
  reg [(5'h11):(1'h0)] reg193 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg192 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg191 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg190 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg189 = (1'h0);
  reg [(5'h10):(1'h0)] forvar222 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg218 = (1'h0);
  reg [(4'ha):(1'h0)] forvar214 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg213 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg212 = (1'h0);
  reg [(5'h13):(1'h0)] reg200 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg194 = (1'h0);
  assign y = {wire225,
                 wire224,
                 wire187,
                 reg223,
                 reg221,
                 reg220,
                 reg219,
                 reg217,
                 reg216,
                 reg215,
                 reg211,
                 reg210,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg199,
                 reg198,
                 reg197,
                 reg196,
                 reg195,
                 reg193,
                 reg192,
                 reg191,
                 reg190,
                 reg189,
                 forvar222,
                 reg218,
                 forvar214,
                 reg213,
                 reg212,
                 reg200,
                 reg194,
                 (1'h0)};
  module5 #() modinst188 (.y(wire187), .wire10(wire2), .wire6(wire3), .wire9(wire1), .clk(clk), .wire7(wire0), .wire8(wire4));
  always
    @(posedge clk) begin
      reg189 <= (wire187[(4'h8):(1'h0)] ?
          "aaWVWMQc5dsQBLBsGNlf" : wire0[(4'he):(4'h9)]);
      if (wire2)
        begin
          reg190 <= $signed($signed($signed({(7'h40), {(8'hae), wire4}})));
          reg191 <= (|(8'had));
          reg192 <= (^~reg191[(1'h0):(1'h0)]);
          reg193 <= $signed(reg192[(1'h1):(1'h1)]);
        end
      else
        begin
          reg194 = (wire2[(3'h6):(1'h0)] >> $unsigned($signed($unsigned((reg190 || reg191)))));
        end
      if ({$unsigned("aroPg2xbN3k9sEWQBe")})
        begin
          reg195 <= $unsigned(reg193[(4'h9):(2'h3)]);
          if (({({(8'ha1),
                  wire0[(5'h11):(5'h11)]} + wire3)} <<< (reg190[(1'h0):(1'h0)] ?
              $signed((((8'hab) * wire3) - (^(8'h9d)))) : (8'hae))))
            begin
              reg196 <= "oeGbEF4c4rZMb9g";
            end
          else
            begin
              reg196 <= $signed(($signed({((8'ha9) ? (8'h9f) : (8'hb4)),
                  $signed(wire4)}) >> "hwQQgR4Ot6RYLdtH"));
            end
          reg197 <= ((8'ha0) <<< $unsigned(wire3));
          reg198 <= reg192[(1'h0):(1'h0)];
          reg199 <= {reg196[(3'h6):(2'h3)],
              {wire1, (!{$signed(wire0), (~^reg196)})}};
        end
      else
        begin
          reg195 <= (wire2[(4'hd):(1'h0)] ?
              ((^~"gpCOhRToMQkpQ") >>> ({reg192[(3'h5):(2'h3)],
                  "dri8rB"} != $signed({reg191,
                  (7'h42)}))) : $unsigned((8'haf)));
          reg196 <= reg194;
          reg200 = $unsigned(wire4[(4'h8):(4'h8)]);
        end
      reg201 <= wire187;
    end
  always
    @(posedge clk) begin
      reg202 <= wire0[(3'h4):(2'h3)];
      if (reg197)
        begin
          reg203 <= ($signed((8'hb6)) ?
              reg190[(1'h1):(1'h1)] : {"y5ZSeuXuiJfoXFHMO1fk",
                  (($unsigned((8'hbf)) ?
                      $signed(reg202) : (~|(8'hab))) | {(reg196 | (8'hb6))})});
          reg204 <= {wire1[(4'h9):(4'h8)], reg195[(5'h10):(3'h6)]};
          if (reg195[(3'h5):(2'h2)])
            begin
              reg205 <= "N2CvCCr";
            end
          else
            begin
              reg205 <= (~|((~reg189) ?
                  $signed(((reg199 ?
                      reg193 : reg191) ^~ "EPvwA5w2dK")) : "ZPxVmu0HS5B9K6Z0zJK"));
              reg206 <= $signed("a5z");
              reg207 <= reg206[(4'hb):(4'hb)];
              reg208 <= $signed((-"vnexySm"));
              reg209 <= ($signed((8'hb1)) ?
                  reg207 : ((8'hb6) ?
                      $signed("Uvum9DDZh15pTJhE") : (($unsigned((8'had)) == reg190) ?
                          (8'h9e) : "t2RTX")));
            end
          reg210 <= ($signed((~|((8'hbd) & $unsigned((8'hb6))))) > "dUHu");
          reg211 <= (~^"cEFJ9SWNwmmD");
        end
      else
        begin
          reg203 <= (reg202[(5'h11):(2'h2)] ~^ $signed(((((8'h9f) ?
                  reg201 : (8'haf)) ?
              $unsigned((8'ha5)) : (7'h41)) - $signed((|(8'hb2))))));
          reg204 <= (^{{(reg196[(5'h11):(4'ha)] ? (8'ha5) : reg204)}, (8'had)});
          reg212 = {$unsigned({reg197[(2'h2):(2'h2)]})};
          reg213 = "oZHZug";
          for (forvar214 = (1'h0); (forvar214 < (2'h2)); forvar214 = (forvar214 + (1'h1)))
            begin
              reg215 <= "y4w6dhlUSibiCLA";
              reg216 <= $unsigned($unsigned(reg205));
              reg217 <= reg204[(1'h0):(1'h0)];
              reg218 = reg191;
              reg219 <= (|reg201);
            end
        end
      reg220 <= $signed(({$unsigned((^~reg216))} ^~ ($unsigned((&(8'ha6))) != reg206[(4'ha):(2'h2)])));
      reg221 <= $signed(reg189[(4'hf):(2'h2)]);
      for (forvar222 = (1'h0); (forvar222 < (2'h2)); forvar222 = (forvar222 + (1'h1)))
        begin
          reg223 <= $signed((8'ha2));
        end
    end
  assign wire224 = (~|(8'hb7));
  assign wire225 = (wire4[(3'h5):(2'h2)] ?
                       reg211[(2'h3):(2'h3)] : (-wire1[(4'hb):(4'hb)]));
endmodule

module module5
#(parameter param185 = (8'hba), 
parameter param186 = ((~({(8'hb9), {(7'h43), param185}} || param185)) <<< param185))
(y, clk, wire6, wire7, wire8, wire9, wire10);
  output wire [(32'h47):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire6;
  input wire [(4'h9):(1'h0)] wire7;
  input wire [(3'h5):(1'h0)] wire8;
  input wire signed [(4'hd):(1'h0)] wire9;
  input wire [(5'h12):(1'h0)] wire10;
  wire signed [(4'ha):(1'h0)] wire184;
  wire signed [(4'hd):(1'h0)] wire183;
  wire signed [(4'hf):(1'h0)] wire182;
  wire [(2'h3):(1'h0)] wire180;
  wire signed [(5'h15):(1'h0)] wire71;
  wire signed [(4'h8):(1'h0)] wire69;
  assign y = {wire184, wire183, wire182, wire180, wire71, wire69, (1'h0)};
  module11 #() modinst70 (.y(wire69), .clk(clk), .wire16(wire9), .wire12(wire8), .wire13(wire10), .wire14(wire7), .wire15(wire6));
  assign wire71 = (!$signed($unsigned($signed("tkzLuM"))));
  module72 #() modinst181 (.wire75(wire10), .wire73(wire8), .wire76(wire71), .clk(clk), .y(wire180), .wire74(wire69));
  assign wire182 = "";
  assign wire183 = wire71;
  assign wire184 = {$unsigned($unsigned((^wire180)))};
endmodule

module module72  (y, clk, wire76, wire75, wire74, wire73);
  output wire [(32'h514):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h4):(1'h0)] wire76;
  input wire [(5'h12):(1'h0)] wire75;
  input wire [(3'h4):(1'h0)] wire74;
  input wire [(3'h5):(1'h0)] wire73;
  wire signed [(3'h7):(1'h0)] wire179;
  wire signed [(4'he):(1'h0)] wire171;
  wire [(5'h12):(1'h0)] wire144;
  wire signed [(4'hb):(1'h0)] wire104;
  wire [(5'h15):(1'h0)] wire91;
  reg signed [(5'h15):(1'h0)] reg178 = (1'h0);
  reg [(5'h13):(1'h0)] reg176 = (1'h0);
  reg [(3'h4):(1'h0)] reg175 = (1'h0);
  reg [(4'hb):(1'h0)] reg174 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg170 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg169 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg168 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg167 = (1'h0);
  reg [(4'h9):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg163 = (1'h0);
  reg [(4'hd):(1'h0)] reg162 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg161 = (1'h0);
  reg [(2'h2):(1'h0)] reg160 = (1'h0);
  reg [(4'he):(1'h0)] reg159 = (1'h0);
  reg [(5'h12):(1'h0)] reg158 = (1'h0);
  reg [(4'hc):(1'h0)] reg157 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg155 = (1'h0);
  reg [(3'h7):(1'h0)] reg153 = (1'h0);
  reg [(4'h9):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg150 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg149 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg146 = (1'h0);
  reg [(5'h10):(1'h0)] reg145 = (1'h0);
  reg [(5'h14):(1'h0)] reg143 = (1'h0);
  reg [(4'hf):(1'h0)] reg142 = (1'h0);
  reg [(5'h15):(1'h0)] reg140 = (1'h0);
  reg [(4'he):(1'h0)] reg138 = (1'h0);
  reg [(4'hf):(1'h0)] reg136 = (1'h0);
  reg signed [(4'he):(1'h0)] reg135 = (1'h0);
  reg [(2'h3):(1'h0)] reg134 = (1'h0);
  reg [(5'h13):(1'h0)] reg133 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg132 = (1'h0);
  reg [(5'h11):(1'h0)] reg129 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg128 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg127 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg126 = (1'h0);
  reg [(3'h7):(1'h0)] reg125 = (1'h0);
  reg [(5'h13):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg121 = (1'h0);
  reg [(5'h12):(1'h0)] reg120 = (1'h0);
  reg [(4'hc):(1'h0)] reg119 = (1'h0);
  reg [(4'ha):(1'h0)] reg118 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg116 = (1'h0);
  reg [(5'h15):(1'h0)] reg115 = (1'h0);
  reg [(5'h11):(1'h0)] reg114 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg111 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg110 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg108 = (1'h0);
  reg [(5'h10):(1'h0)] reg105 = (1'h0);
  reg [(5'h15):(1'h0)] reg102 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg101 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg100 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg98 = (1'h0);
  reg [(3'h7):(1'h0)] reg97 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg96 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg95 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg94 = (1'h0);
  reg [(4'hd):(1'h0)] reg93 = (1'h0);
  reg [(4'hf):(1'h0)] reg92 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg90 = (1'h0);
  reg [(4'hc):(1'h0)] reg89 = (1'h0);
  reg [(4'hd):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg87 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg84 = (1'h0);
  reg [(4'hd):(1'h0)] reg77 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg82 = (1'h0);
  reg [(2'h2):(1'h0)] reg81 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg80 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg79 = (1'h0);
  reg [(2'h3):(1'h0)] reg78 = (1'h0);
  reg [(3'h4):(1'h0)] reg177 = (1'h0);
  reg [(4'hb):(1'h0)] forvar173 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar172 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg166 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar165 = (1'h0);
  reg [(2'h3):(1'h0)] reg156 = (1'h0);
  reg [(5'h11):(1'h0)] forvar154 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg152 = (1'h0);
  reg [(4'ha):(1'h0)] reg148 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg147 = (1'h0);
  reg [(4'hf):(1'h0)] reg141 = (1'h0);
  reg [(4'hf):(1'h0)] forvar139 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg137 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar131 = (1'h0);
  reg [(3'h5):(1'h0)] forvar130 = (1'h0);
  reg [(5'h11):(1'h0)] reg124 = (1'h0);
  reg [(3'h5):(1'h0)] forvar123 = (1'h0);
  reg [(4'hc):(1'h0)] reg122 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar117 = (1'h0);
  reg [(4'hf):(1'h0)] reg112 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar106 = (1'h0);
  reg [(2'h2):(1'h0)] reg103 = (1'h0);
  reg [(5'h14):(1'h0)] forvar99 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg86 = (1'h0);
  reg [(2'h3):(1'h0)] forvar85 = (1'h0);
  reg [(3'h5):(1'h0)] reg83 = (1'h0);
  reg [(4'ha):(1'h0)] forvar77 = (1'h0);
  assign y = {wire179,
                 wire171,
                 wire144,
                 wire104,
                 wire91,
                 reg178,
                 reg176,
                 reg175,
                 reg174,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg164,
                 reg163,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg158,
                 reg157,
                 reg155,
                 reg153,
                 reg151,
                 reg150,
                 reg149,
                 reg146,
                 reg145,
                 reg143,
                 reg142,
                 reg140,
                 reg138,
                 reg136,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg129,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg123,
                 reg121,
                 reg120,
                 reg119,
                 reg118,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg105,
                 reg102,
                 reg101,
                 reg100,
                 reg98,
                 reg97,
                 reg96,
                 reg95,
                 reg94,
                 reg93,
                 reg92,
                 reg90,
                 reg89,
                 reg88,
                 reg87,
                 reg84,
                 reg77,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg78,
                 reg177,
                 forvar173,
                 forvar172,
                 reg166,
                 forvar165,
                 reg156,
                 forvar154,
                 reg152,
                 reg148,
                 reg147,
                 reg141,
                 forvar139,
                 reg137,
                 forvar131,
                 forvar130,
                 reg124,
                 forvar123,
                 reg122,
                 forvar117,
                 reg112,
                 reg107,
                 forvar106,
                 reg103,
                 forvar99,
                 reg86,
                 forvar85,
                 reg83,
                 forvar77,
                 (1'h0)};
  always
    @(posedge clk) begin
      if (wire73)
        begin
          for (forvar77 = (1'h0); (forvar77 < (3'h4)); forvar77 = (forvar77 + (1'h1)))
            begin
              reg78 <= $unsigned($unsigned("SpxFZiPsZq6xPlU1x"));
            end
          reg79 <= wire74[(1'h1):(1'h0)];
          if ((~^{(8'ha7),
              (($signed(wire76) ? reg78 : (~&wire75)) ?
                  forvar77 : ({(8'hac)} ? "bZVUJ" : (wire73 << wire75)))}))
            begin
              reg80 <= $signed((wire76 ? (^~(8'hab)) : $signed(wire74)));
              reg81 <= reg80[(4'ha):(3'h4)];
              reg82 <= $signed($unsigned(((7'h43) ?
                  (reg80 << (|reg79)) : (8'had))));
            end
          else
            begin
              reg80 <= $unsigned(forvar77[(1'h1):(1'h0)]);
              reg81 <= ((8'h9c) >= reg80[(4'h8):(3'h5)]);
            end
          reg83 = ({(+reg82[(4'ha):(1'h1)]),
                  ($signed(wire76[(3'h4):(2'h2)]) ?
                      $unsigned(((8'hb5) ? wire74 : (8'h9f))) : ((7'h43) ?
                          "urM3ZYH0fwEs" : {(8'hb6), (8'ha4)}))} ?
              wire73[(2'h2):(1'h1)] : forvar77);
        end
      else
        begin
          reg77 <= $unsigned((8'ha4));
          reg78 <= "3zGLJ7P0l7hN0W3inW";
          reg83 = (&(($signed({wire76, wire74}) < ({wire76} ?
                  ((8'hb4) << (8'hb7)) : $signed(reg82))) ?
              $unsigned(("aZdMnI" ^~ wire73[(3'h5):(3'h5)])) : {reg79[(2'h2):(1'h1)],
                  (+(reg82 && reg80))}));
        end
      reg84 <= "JwAYXvQL0564";
      for (forvar85 = (1'h0); (forvar85 < (1'h1)); forvar85 = (forvar85 + (1'h1)))
        begin
          reg86 = (($unsigned($unsigned($unsigned((8'h9e)))) || reg81) >> "hXKJo5azTG");
          reg87 <= (($unsigned($unsigned((reg79 <= reg79))) ?
              (wire73 | ({reg77, (8'h9f)} ?
                  (8'hbb) : reg83[(1'h0):(1'h0)])) : (8'ha8)) ^~ "sfpIx");
          reg88 <= (^(((!{(8'h9f)}) ? "2" : $signed(((8'hb3) << (8'hbc)))) ?
              (8'ha0) : "rzbQQlWJEB"));
        end
      reg89 <= $signed((wire73[(3'h4):(1'h0)] * "bSiobJpYgGQu"));
      reg90 <= $signed(reg86[(5'h13):(4'hd)]);
    end
  assign wire91 = $signed(("3w" ?
                      reg78[(2'h3):(1'h1)] : ((^~(8'hb9)) ?
                          "" : (reg78 ?
                              ((8'hb6) ? (8'ha2) : (8'hab)) : (^reg78)))));
  always
    @(posedge clk) begin
      reg92 <= $unsigned($unsigned((8'ha1)));
      reg93 <= (~$unsigned((&(wire91 ?
          ((8'ha2) ? reg84 : (8'ha7)) : "Ep25r"))));
      reg94 <= "19ipo";
      if (reg92[(2'h2):(1'h1)])
        begin
          reg95 <= wire75[(3'h5):(1'h0)];
          reg96 <= $signed($unsigned(wire76));
        end
      else
        begin
          reg95 <= $signed($signed((8'haa)));
        end
      reg97 <= (+$unsigned($unsigned(((wire76 <= (8'hb0)) ?
          (8'hae) : "gWzY1Y1"))));
    end
  always
    @(posedge clk) begin
      reg98 <= (8'hba);
      for (forvar99 = (1'h0); (forvar99 < (3'h4)); forvar99 = (forvar99 + (1'h1)))
        begin
          reg100 <= "RvwCoOtwIZdqa3J46";
          reg101 <= $unsigned($unsigned(reg84[(1'h0):(1'h0)]));
        end
      reg102 <= $unsigned((8'hb2));
      reg103 = {(("xYkJtlrphkBEeXz" ?
                  $unsigned((reg78 ? wire75 : (8'haf))) : {"CDPbUJcRHsGXDxt",
                      (reg95 < reg92)}) ?
              ({((8'hb4) ? (8'hb0) : reg84)} << (7'h42)) : $unsigned({wire75,
                  (~&(8'ha7))})),
          (reg93[(2'h3):(2'h2)] ?
              "VZLfCM" : (($unsigned(reg94) - ((7'h44) ? (8'hb1) : (8'hb7))) ?
                  wire91 : (8'h9c)))};
    end
  assign wire104 = (8'hab);
  always
    @(posedge clk) begin
      reg105 <= (8'hbf);
    end
  always
    @(posedge clk) begin
      for (forvar106 = (1'h0); (forvar106 < (2'h2)); forvar106 = (forvar106 + (1'h1)))
        begin
          reg107 = reg81[(1'h1):(1'h0)];
          reg108 <= wire74[(2'h3):(2'h3)];
          if ((({(8'ha3)} ? "rfGvD4GUXV" : $signed($signed({wire76}))) ^~ ""))
            begin
              reg109 <= "1Ivt";
              reg110 <= {reg101, (8'ha8)};
              reg111 <= "NLD2RdAgaL3hAb59";
            end
          else
            begin
              reg112 = reg78[(2'h2):(1'h1)];
              reg113 <= $unsigned((reg89[(3'h5):(2'h3)] || "PLIS"));
              reg114 <= $unsigned(reg102[(3'h4):(3'h4)]);
              reg115 <= ((8'hac) == $signed(("gKP" ^~ $signed((8'hbc)))));
            end
        end
      reg116 <= (reg95 ?
          ((8'hbf) * (^~(^wire73))) : $unsigned(reg97[(3'h5):(2'h3)]));
      for (forvar117 = (1'h0); (forvar117 < (2'h3)); forvar117 = (forvar117 + (1'h1)))
        begin
          reg118 <= ((&reg113) && (8'hb1));
          reg119 <= reg111[(1'h0):(1'h0)];
          reg120 <= (reg77 ? ("0D3" | forvar106) : reg119);
          reg121 <= $unsigned((+(7'h41)));
        end
      reg122 = {(reg105 ?
              $signed((|$signed(forvar106))) : reg101[(4'h9):(4'h8)]),
          {(7'h42), (^reg77)}};
    end
  always
    @(posedge clk) begin
      if (($signed(reg105) ? reg87 : reg114[(5'h10):(4'hc)]))
        begin
          for (forvar123 = (1'h0); (forvar123 < (1'h0)); forvar123 = (forvar123 + (1'h1)))
            begin
              reg124 = (8'hb0);
            end
        end
      else
        begin
          reg123 <= (wire76[(2'h2):(2'h2)] ?
              (((^~(~^reg116)) ?
                  reg114[(4'ha):(4'h8)] : ((~|reg78) ?
                      (-reg78) : {reg113})) * (-"sLwzpaRDkU")) : ((!(8'hb0)) ?
                  ("HNkqh9b3NqD" ?
                      (^~wire75) : "hovnBtpsKdanNwu") : $signed(($signed((8'hac)) ?
                      (8'ha4) : ((8'ha8) << reg97)))));
          reg125 <= (8'hb6);
          reg126 <= $signed($signed((8'hb2)));
          reg127 <= reg88;
          reg128 <= ($signed(reg108[(4'hf):(4'he)]) ?
              {(reg110[(1'h1):(1'h0)] ?
                      ($signed((8'ha3)) ?
                          wire104 : ((8'ha8) ?
                              (8'hbd) : reg113)) : (reg92 == {(8'hbc),
                          (8'ha2)})),
                  reg80} : ((7'h44) & wire75));
        end
      reg129 <= ((8'haa) ~^ (8'ha6));
      for (forvar130 = (1'h0); (forvar130 < (2'h3)); forvar130 = (forvar130 + (1'h1)))
        begin
          for (forvar131 = (1'h0); (forvar131 < (3'h4)); forvar131 = (forvar131 + (1'h1)))
            begin
              reg132 <= $unsigned((8'ha9));
              reg133 <= $unsigned(reg87[(4'hc):(1'h1)]);
              reg134 <= wire76[(2'h2):(2'h2)];
              reg135 <= (~^{(8'ha8), (8'hb8)});
              reg136 <= $unsigned((($unsigned($unsigned((8'ha5))) != $signed($signed((8'hae)))) >> $unsigned(((reg127 ^~ reg89) * $signed(reg116)))));
            end
          reg137 = $signed((8'h9e));
          reg138 <= (((8'hae) << $signed((!(reg94 ?
              (8'ha5) : reg123)))) + (^~"DgMXp9RzI"));
          for (forvar139 = (1'h0); (forvar139 < (3'h4)); forvar139 = (forvar139 + (1'h1)))
            begin
              reg140 <= $signed(reg94[(2'h3):(2'h3)]);
              reg141 = ($signed((~|$unsigned(reg90))) ?
                  reg133[(4'hf):(1'h1)] : reg82);
              reg142 <= reg101[(3'h7):(3'h6)];
            end
        end
      reg143 <= "lr64RSTFiNfo6";
    end
  assign wire144 = ((-"iwfo2CX") ? "HprnCKi32s04HBaz6zr" : $unsigned(reg80));
  always
    @(posedge clk) begin
      reg145 <= ("XV9Ee5mbkP7xGid08lZF" > wire74[(2'h3):(2'h3)]);
      reg146 <= (8'ha5);
      reg147 = (^$signed(wire144[(4'hf):(4'hb)]));
    end
  always
    @(posedge clk) begin
      reg148 = wire91;
      reg149 <= $unsigned(reg97[(3'h5):(3'h5)]);
      reg150 <= reg119;
      reg151 <= reg127;
      reg152 = wire76[(2'h2):(1'h1)];
    end
  always
    @(posedge clk) begin
      reg153 <= $unsigned($signed((reg128 ^~ wire74[(2'h2):(1'h1)])));
      for (forvar154 = (1'h0); (forvar154 < (2'h2)); forvar154 = (forvar154 + (1'h1)))
        begin
          if (reg84[(1'h0):(1'h0)])
            begin
              reg155 <= (!(~^{({reg134} >>> reg113),
                  ({reg95} | "6t45NEAboeZ8")}));
              reg156 = {($unsigned($unsigned((8'hb2))) ?
                      (7'h40) : "smhstLyIEnMgutoes"),
                  (^((reg119 & "Lqebna2L8rhtAt6") & $signed(((8'haf) * (8'hb8)))))};
              reg157 <= {($signed("") <= $signed((^$signed((8'hbf))))), reg81};
              reg158 <= (((7'h42) >= (wire74[(2'h3):(2'h3)] < $signed(reg95))) ?
                  ((reg102[(5'h13):(3'h4)] ?
                          {reg80[(1'h0):(1'h0)]} : (((8'hab) + (8'hae)) ?
                              $unsigned((8'hbd)) : reg92)) ?
                      "65sp4QzRS0Mr1C" : "ZkMbO") : reg88);
            end
          else
            begin
              reg156 = "upKUgPRcWyxny56N";
              reg157 <= (|reg102[(2'h2):(1'h0)]);
              reg158 <= {$signed((-(^~(reg157 >>> reg121)))),
                  reg129[(3'h4):(1'h1)]};
              reg159 <= (!(((!"mbSpGdyFMg23") | ((reg114 << reg93) ?
                      (|reg129) : (~&wire76))) ?
                  $signed(reg142[(1'h0):(1'h0)]) : (~^(~$unsigned((8'hb8))))));
              reg160 <= $signed(reg87);
            end
          if ($signed((($unsigned((reg136 < reg129)) >= (!((8'hae) >> reg108))) ?
              ({$unsigned(reg110)} ?
                  (reg151[(2'h3):(1'h1)] | (8'ha5)) : (~|$unsigned((8'ha3)))) : (|(+reg155)))))
            begin
              reg161 <= reg127[(3'h6):(1'h1)];
              reg162 <= ($signed(($signed((reg108 ?
                      reg90 : (8'hb0))) >> reg160)) ?
                  (((reg88 << reg156[(1'h0):(1'h0)]) << (!$signed((8'hab)))) ?
                      "F6s9CKLsx4" : (reg100[(2'h2):(1'h0)] ?
                          wire104[(4'h9):(3'h5)] : ("pWZr1du2S" + (~(8'ha7))))) : (wire91[(5'h12):(1'h1)] ^ ((8'ha5) ?
                      $unsigned(reg129[(4'he):(1'h1)]) : (^reg160))));
              reg163 <= reg95[(5'h11):(4'hf)];
              reg164 <= $signed($signed(($signed((reg92 != (7'h44))) ?
                  {reg149} : reg108)));
            end
          else
            begin
              reg161 <= (wire104[(4'h9):(4'h8)] ? reg125 : reg159);
            end
          for (forvar165 = (1'h0); (forvar165 < (2'h3)); forvar165 = (forvar165 + (1'h1)))
            begin
              reg166 = (~&(8'hb1));
              reg167 <= ($signed("ain7qcJi") ?
                  $signed((-$signed("NGBCT2xBr9O32fUg"))) : reg79[(3'h6):(3'h6)]);
              reg168 <= ($signed({reg160,
                  "26SMK5JrXC"}) >= $signed(reg77[(1'h0):(1'h0)]));
            end
        end
      reg169 <= $signed(((8'hae) ?
          {(((8'hb7) ^~ reg127) >> (reg82 || (8'h9f)))} : (reg119 >> {((8'ha8) ?
                  reg149 : (8'ha0))})));
    end
  always
    @(posedge clk) begin
      reg170 <= reg78;
    end
  assign wire171 = $signed($signed(reg84[(2'h2):(2'h2)]));
  always
    @(posedge clk) begin
      for (forvar172 = (1'h0); (forvar172 < (2'h2)); forvar172 = (forvar172 + (1'h1)))
        begin
          for (forvar173 = (1'h0); (forvar173 < (1'h0)); forvar173 = (forvar173 + (1'h1)))
            begin
              reg174 <= reg153;
              reg175 <= reg92[(4'hb):(2'h2)];
              reg176 <= ((~&((8'hb1) != $signed($signed(reg88)))) & (("6bb8R" == ("ZlGhPwpmfY0N" || (8'ha4))) ?
                  (~|(8'haa)) : (~^(~^wire75[(3'h5):(1'h1)]))));
              reg177 = $unsigned($unsigned(reg136));
              reg178 <= (|(8'ha3));
            end
        end
    end
  assign wire179 = "sD7F0";
endmodule

module module11
#(parameter param68 = ((((8'haf) >> ((-(8'hb3)) ? (8'hba) : ((8'h9e) ? (7'h40) : (8'hb8)))) | (8'ha0)) ? (8'ha0) : (~&(8'ha0))))
(y, clk, wire16, wire15, wire14, wire13, wire12);
  output wire [(32'h23f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h3):(1'h0)] wire16;
  input wire signed [(4'hb):(1'h0)] wire15;
  input wire [(2'h3):(1'h0)] wire14;
  input wire signed [(3'h5):(1'h0)] wire13;
  input wire [(2'h3):(1'h0)] wire12;
  wire signed [(5'h14):(1'h0)] wire49;
  wire signed [(5'h12):(1'h0)] wire17;
  reg [(4'hc):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg66 = (1'h0);
  reg [(3'h7):(1'h0)] reg65 = (1'h0);
  reg [(3'h4):(1'h0)] reg64 = (1'h0);
  reg [(5'h14):(1'h0)] reg63 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg62 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg61 = (1'h0);
  reg [(5'h10):(1'h0)] reg58 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg56 = (1'h0);
  reg [(5'h11):(1'h0)] reg54 = (1'h0);
  reg [(4'h9):(1'h0)] reg53 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg52 = (1'h0);
  reg [(2'h3):(1'h0)] reg48 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg44 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg43 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg41 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg40 = (1'h0);
  reg [(4'h8):(1'h0)] reg38 = (1'h0);
  reg [(2'h2):(1'h0)] reg36 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg35 = (1'h0);
  reg [(4'hc):(1'h0)] reg34 = (1'h0);
  reg [(5'h14):(1'h0)] reg33 = (1'h0);
  reg [(5'h14):(1'h0)] reg32 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg31 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg30 = (1'h0);
  reg [(2'h3):(1'h0)] reg29 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg28 = (1'h0);
  reg [(5'h10):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg26 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg24 = (1'h0);
  reg [(5'h15):(1'h0)] reg23 = (1'h0);
  reg [(5'h15):(1'h0)] reg21 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg20 = (1'h0);
  reg [(5'h15):(1'h0)] reg18 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar60 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg59 = (1'h0);
  reg [(5'h11):(1'h0)] reg55 = (1'h0);
  reg [(4'hf):(1'h0)] reg51 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar50 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg47 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg46 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg45 = (1'h0);
  reg [(4'h9):(1'h0)] forvar42 = (1'h0);
  reg [(3'h5):(1'h0)] reg39 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg37 = (1'h0);
  reg [(2'h2):(1'h0)] reg25 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar22 = (1'h0);
  reg [(4'h9):(1'h0)] forvar19 = (1'h0);
  assign y = {wire49,
                 wire17,
                 reg67,
                 reg66,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg61,
                 reg58,
                 reg57,
                 reg56,
                 reg54,
                 reg53,
                 reg52,
                 reg48,
                 reg44,
                 reg43,
                 reg41,
                 reg40,
                 reg38,
                 reg36,
                 reg35,
                 reg34,
                 reg33,
                 reg32,
                 reg31,
                 reg30,
                 reg29,
                 reg28,
                 reg27,
                 reg26,
                 reg24,
                 reg23,
                 reg21,
                 reg20,
                 reg18,
                 forvar60,
                 reg59,
                 reg55,
                 reg51,
                 forvar50,
                 reg47,
                 reg46,
                 reg45,
                 forvar42,
                 reg39,
                 reg37,
                 reg25,
                 forvar22,
                 forvar19,
                 (1'h0)};
  assign wire17 = (wire14[(1'h0):(1'h0)] ^~ $signed(wire15[(4'ha):(3'h6)]));
  always
    @(posedge clk) begin
      reg18 <= "qmHZUAr5HV9cMWLO";
      for (forvar19 = (1'h0); (forvar19 < (1'h0)); forvar19 = (forvar19 + (1'h1)))
        begin
          reg20 <= $signed((wire13 ?
              "tK7wa9tun8JqQDR" : ((8'ha6) ?
                  $signed($signed((8'haa))) : ({(8'ha1), wire17} != (8'ha6)))));
          reg21 <= ({((8'hb5) ? (|(8'hb8)) : (forvar19 ? "aBMI1Dde6FWP" : "Z")),
                  (8'hb1)} ?
              (((+((8'ha4) ? wire13 : reg18)) ?
                  $signed(reg18) : $unsigned($unsigned((8'ha6)))) * (8'h9d)) : wire14);
          for (forvar22 = (1'h0); (forvar22 < (2'h2)); forvar22 = (forvar22 + (1'h1)))
            begin
              reg23 <= $unsigned(((wire13[(3'h4):(1'h1)] >>> $signed($unsigned((8'hb6)))) ?
                  (~|wire16[(1'h1):(1'h0)]) : (~|($signed(wire16) ^~ $unsigned((8'ha0))))));
              reg24 <= ($unsigned((8'hbf)) >= (8'h9e));
            end
          reg25 = (8'ha3);
        end
      reg26 <= (($signed(wire17) < $unsigned((^(wire12 - (8'had))))) != (wire14[(2'h3):(2'h3)] ?
          $unsigned(wire16[(2'h3):(2'h2)]) : $signed(reg18[(3'h6):(3'h4)])));
      reg27 <= reg25;
    end
  always
    @(posedge clk) begin
      reg28 <= $signed(((~|(wire16 ?
          reg24 : $signed(reg27))) == wire15[(3'h7):(3'h6)]));
      if ($unsigned({((&(|reg26)) + $unsigned(reg21[(3'h5):(3'h5)])),
          (reg26[(5'h10):(4'hf)] ? (8'haf) : $signed(((8'hb3) ^~ (8'hb0))))}))
        begin
          reg29 <= "fVXxf8doNV48VDu";
          reg30 <= "mWU";
          reg31 <= $unsigned(wire13);
        end
      else
        begin
          reg29 <= "";
          reg30 <= (8'ha2);
        end
      reg32 <= ((($unsigned($signed((8'hbe))) << $unsigned(wire16)) >> wire15) <<< $unsigned(reg21[(4'h9):(3'h5)]));
      reg33 <= (7'h42);
      reg34 <= "4K8I";
    end
  always
    @(posedge clk) begin
      reg35 <= (((^{"ASfyKE5ctBJ9", reg28}) * (8'hb2)) - ((8'hb3) ?
          reg20[(3'h5):(1'h0)] : reg18[(5'h10):(4'hf)]));
      reg36 <= "ydh5J8ctXWf";
      if (($signed((reg35[(1'h1):(1'h0)] & wire16)) >> ((reg35[(1'h1):(1'h1)] >= reg29) - "sNGQ2")))
        begin
          reg37 = (~|$signed(((8'hb3) ?
              (7'h40) : (((8'h9f) >= (8'hbe)) ? reg23 : $unsigned((8'h9d))))));
          reg38 <= $unsigned((~(7'h40)));
        end
      else
        begin
          reg38 <= reg24[(3'h7):(3'h7)];
          reg39 = $unsigned(((reg26[(4'h9):(3'h6)] ?
                  "QX6RoIP" : (^~reg36[(1'h0):(1'h0)])) ?
              $signed(($unsigned(reg30) ?
                  "9WY" : ((8'hbf) ? (8'ha9) : (8'hb6)))) : reg27));
          reg40 <= ((~^{(8'ha3), "Nzrb"}) ?
              ("SdtOmYVbGLdl5UlCQ6" ?
                  wire12 : $unsigned(((reg29 ? reg39 : (8'hb0)) ?
                      reg32 : ((8'hb6) && wire13)))) : ((reg18[(4'hb):(2'h3)] ?
                      ((~^reg20) ?
                          $signed((8'ha2)) : reg33[(2'h2):(2'h2)]) : "D") ?
                  (8'h9f) : {wire14[(2'h2):(1'h1)]}));
        end
      reg41 <= $unsigned(reg34[(4'h8):(2'h3)]);
      if ($unsigned({(((~^(8'hb4)) ? reg24 : reg39) - $unsigned("")),
          "L7Srf9k0ruAXZT97XqAe"}))
        begin
          for (forvar42 = (1'h0); (forvar42 < (2'h2)); forvar42 = (forvar42 + (1'h1)))
            begin
              reg43 <= "5QNAYbnBRLBGcAeVlQfP";
              reg44 <= $signed($signed(((8'ha1) >= ($signed((8'ha8)) | reg40[(3'h4):(2'h2)]))));
            end
          reg45 = (({reg35} ?
                  ("7aJ4SsGPfisPreL" ?
                      ((+(8'hb9)) >= ((7'h41) ? wire15 : (8'ha7))) : (((7'h44) ?
                              (8'had) : reg37) ?
                          $unsigned(reg35) : (&reg24))) : $unsigned(reg37)) ?
              $signed($unsigned({((8'hac) ? (8'hae) : wire12),
                  $unsigned((8'haa))})) : $unsigned((reg38 >> (8'h9e))));
          reg46 = (reg29 ? (8'hb9) : $signed(wire17[(1'h0):(1'h0)]));
          reg47 = $unsigned(reg24[(2'h2):(1'h0)]);
        end
      else
        begin
          for (forvar42 = (1'h0); (forvar42 < (2'h2)); forvar42 = (forvar42 + (1'h1)))
            begin
              reg43 <= wire12[(2'h2):(1'h1)];
              reg44 <= (8'hb9);
              reg45 = {$unsigned(("INBKIgLyuzu4FzV" ?
                      {(~(8'h9f))} : forvar42))};
            end
          reg48 <= (8'hbe);
        end
    end
  assign wire49 = reg44[(3'h4):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar50 = (1'h0); (forvar50 < (2'h3)); forvar50 = (forvar50 + (1'h1)))
        begin
          if (wire17)
            begin
              reg51 = ((($signed(((8'hb6) + reg18)) ?
                      ($signed(wire12) >>> $signed(reg23)) : (wire17 != forvar50)) > reg26) ?
                  "wTcCoPGIWAy" : (8'ha2));
            end
          else
            begin
              reg52 <= ((reg32[(3'h4):(1'h1)] ?
                      (((reg48 ? reg35 : wire15) ?
                          wire15[(4'h8):(3'h5)] : (8'haa)) != (8'hb8)) : (reg21 || ((reg28 ?
                              (8'hb7) : reg48) ?
                          $signed((8'ha4)) : (8'hba)))) ?
                  (8'ha4) : "GL7aIb7OV56ZWVKEGd");
              reg53 <= reg30;
              reg54 <= wire17[(4'h9):(3'h4)];
              reg55 = "u6cMA0nzpnSTb2Fpu";
            end
          reg56 <= (reg28 ? (7'h40) : reg28[(3'h5):(2'h3)]);
          reg57 <= (~^((~&reg38) >> ((&((8'hb4) + (7'h43))) > $unsigned((~|(8'hb4))))));
          reg58 <= $signed({reg48});
          reg59 = (~^(~^wire15[(3'h5):(3'h5)]));
        end
      for (forvar60 = (1'h0); (forvar60 < (2'h3)); forvar60 = (forvar60 + (1'h1)))
        begin
          reg61 <= {reg40};
          reg62 <= "r7";
          reg63 <= $unsigned($signed(((8'hb4) >= ((reg43 ?
              wire13 : (8'h9d)) & reg61[(3'h5):(2'h2)]))));
          reg64 <= reg52[(1'h1):(1'h1)];
        end
      reg65 <= reg29[(2'h2):(1'h1)];
      reg66 <= (reg48[(2'h2):(2'h2)] ^~ (reg33 || ("BnkyJczDpxzQycIzReq" != {(!reg24)})));
    end
  always
    @(posedge clk) begin
      reg67 <= (($unsigned("pHfzTU4QHTnrXqqa") ?
          (~^(8'hac)) : $unsigned(reg34)) ~^ reg38);
    end
endmodule