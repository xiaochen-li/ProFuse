(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param607 = {(8'hab)}, 
parameter param608 = (param607 ? ((((param607 ^ param607) > {param607, param607}) & param607) ? (~|(((8'hb5) ? param607 : param607) ? {param607} : param607)) : param607) : (param607 <<< {param607, param607})))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'h565):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire3;
  input wire [(5'h12):(1'h0)] wire2;
  input wire [(4'hf):(1'h0)] wire1;
  input wire [(4'h9):(1'h0)] wire0;
  wire [(2'h2):(1'h0)] wire559;
  wire [(4'h9):(1'h0)] wire558;
  wire [(5'h14):(1'h0)] wire513;
  wire signed [(4'h9):(1'h0)] wire4;
  wire [(4'hb):(1'h0)] wire515;
  wire [(4'he):(1'h0)] wire517;
  wire signed [(4'ha):(1'h0)] wire519;
  wire [(4'h8):(1'h0)] wire520;
  wire signed [(4'hb):(1'h0)] wire521;
  reg signed [(5'h12):(1'h0)] reg606 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg605 = (1'h0);
  reg [(4'h8):(1'h0)] reg604 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg602 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg601 = (1'h0);
  reg [(4'he):(1'h0)] reg599 = (1'h0);
  reg [(5'h12):(1'h0)] reg598 = (1'h0);
  reg [(2'h3):(1'h0)] reg597 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg596 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg593 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg592 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg591 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg590 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg587 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg586 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg585 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg584 = (1'h0);
  reg [(3'h7):(1'h0)] reg583 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg582 = (1'h0);
  reg [(5'h12):(1'h0)] reg581 = (1'h0);
  reg [(5'h14):(1'h0)] reg578 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg577 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg575 = (1'h0);
  reg [(4'h9):(1'h0)] reg574 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg572 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg571 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg570 = (1'h0);
  reg [(5'h12):(1'h0)] reg569 = (1'h0);
  reg [(2'h3):(1'h0)] reg562 = (1'h0);
  reg [(3'h6):(1'h0)] reg567 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg566 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg564 = (1'h0);
  reg [(4'h8):(1'h0)] reg563 = (1'h0);
  reg [(4'hc):(1'h0)] reg5 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg6 = (1'h0);
  reg [(4'hf):(1'h0)] reg8 = (1'h0);
  reg [(5'h14):(1'h0)] reg10 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg11 = (1'h0);
  reg [(3'h4):(1'h0)] reg12 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg13 = (1'h0);
  reg [(5'h11):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg17 = (1'h0);
  reg [(5'h14):(1'h0)] reg18 = (1'h0);
  reg [(4'hc):(1'h0)] reg19 = (1'h0);
  reg [(4'hf):(1'h0)] reg21 = (1'h0);
  reg [(5'h14):(1'h0)] reg22 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg23 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg523 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg524 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg525 = (1'h0);
  reg [(4'h8):(1'h0)] reg526 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg527 = (1'h0);
  reg [(4'he):(1'h0)] reg528 = (1'h0);
  reg [(4'hf):(1'h0)] reg531 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg532 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg533 = (1'h0);
  reg [(4'hc):(1'h0)] reg535 = (1'h0);
  reg [(4'h8):(1'h0)] reg536 = (1'h0);
  reg [(2'h2):(1'h0)] reg537 = (1'h0);
  reg [(2'h2):(1'h0)] reg538 = (1'h0);
  reg [(3'h5):(1'h0)] reg539 = (1'h0);
  reg [(4'hc):(1'h0)] reg541 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg544 = (1'h0);
  reg [(5'h12):(1'h0)] reg545 = (1'h0);
  reg [(4'ha):(1'h0)] reg546 = (1'h0);
  reg [(3'h6):(1'h0)] reg547 = (1'h0);
  reg [(4'he):(1'h0)] reg548 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg549 = (1'h0);
  reg [(4'hd):(1'h0)] reg551 = (1'h0);
  reg [(3'h6):(1'h0)] reg553 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg554 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg555 = (1'h0);
  reg [(3'h4):(1'h0)] reg556 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg557 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg603 = (1'h0);
  reg [(5'h15):(1'h0)] reg600 = (1'h0);
  reg [(3'h6):(1'h0)] forvar594 = (1'h0);
  reg [(4'hd):(1'h0)] reg589 = (1'h0);
  reg [(4'hd):(1'h0)] forvar588 = (1'h0);
  reg [(4'hc):(1'h0)] forvar580 = (1'h0);
  reg [(5'h10):(1'h0)] reg579 = (1'h0);
  reg [(4'hb):(1'h0)] forvar576 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar573 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg568 = (1'h0);
  reg [(3'h6):(1'h0)] forvar565 = (1'h0);
  reg [(5'h13):(1'h0)] forvar562 = (1'h0);
  reg [(3'h7):(1'h0)] reg561 = (1'h0);
  reg [(5'h14):(1'h0)] reg552 = (1'h0);
  reg [(4'ha):(1'h0)] forvar550 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar543 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg542 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar536 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg540 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg534 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar530 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg529 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar525 = (1'h0);
  reg [(5'h13):(1'h0)] reg20 = (1'h0);
  reg [(5'h14):(1'h0)] reg14 = (1'h0);
  reg [(3'h4):(1'h0)] reg9 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar7 = (1'h0);
  assign y = {wire559,
                 wire558,
                 wire513,
                 wire4,
                 wire515,
                 wire517,
                 wire519,
                 wire520,
                 wire521,
                 reg606,
                 reg605,
                 reg604,
                 reg602,
                 reg601,
                 reg599,
                 reg598,
                 reg597,
                 reg596,
                 reg595,
                 reg593,
                 reg592,
                 reg591,
                 reg590,
                 reg587,
                 reg586,
                 reg585,
                 reg584,
                 reg583,
                 reg582,
                 reg581,
                 reg578,
                 reg577,
                 reg575,
                 reg574,
                 reg572,
                 reg571,
                 reg570,
                 reg569,
                 reg562,
                 reg567,
                 reg566,
                 reg564,
                 reg563,
                 reg5,
                 reg6,
                 reg8,
                 reg10,
                 reg11,
                 reg12,
                 reg13,
                 reg15,
                 reg16,
                 reg17,
                 reg18,
                 reg19,
                 reg21,
                 reg22,
                 reg23,
                 reg523,
                 reg524,
                 reg525,
                 reg526,
                 reg527,
                 reg528,
                 reg531,
                 reg532,
                 reg533,
                 reg535,
                 reg536,
                 reg537,
                 reg538,
                 reg539,
                 reg541,
                 reg544,
                 reg545,
                 reg546,
                 reg547,
                 reg548,
                 reg549,
                 reg551,
                 reg553,
                 reg554,
                 reg555,
                 reg556,
                 reg557,
                 reg603,
                 reg600,
                 forvar594,
                 reg589,
                 forvar588,
                 forvar580,
                 reg579,
                 forvar576,
                 forvar573,
                 reg568,
                 forvar565,
                 forvar562,
                 reg561,
                 reg552,
                 forvar550,
                 forvar543,
                 reg542,
                 forvar536,
                 reg540,
                 reg534,
                 forvar530,
                 reg529,
                 forvar525,
                 reg20,
                 reg14,
                 reg9,
                 forvar7,
                 (1'h0)};
  assign wire4 = $unsigned($signed({$signed({wire0, (8'h9d)})}));
  always
    @(posedge clk) begin
      reg5 <= $unsigned({(~|(wire0 ? {wire3, wire3} : $unsigned(wire0))),
          (7'h42)});
      reg6 <= ({(($signed(wire0) ?
              $unsigned(wire3) : (wire4 ? reg5 : reg5)) ^~ wire0)} != wire2);
      for (forvar7 = (1'h0); (forvar7 < (1'h1)); forvar7 = (forvar7 + (1'h1)))
        begin
          reg8 <= $signed(($signed((-wire3[(4'h8):(3'h7)])) * wire0[(3'h6):(1'h1)]));
          reg9 = ($signed($signed($unsigned($signed(forvar7)))) && $unsigned($signed(($unsigned(reg8) ?
              {wire1} : ((8'ha8) ? (8'hb2) : (8'haa))))));
          if (reg5)
            begin
              reg10 <= wire0[(4'h8):(2'h3)];
              reg11 <= {reg9[(1'h0):(1'h0)]};
              reg12 <= $unsigned((!{$unsigned($signed(forvar7))}));
              reg13 <= $unsigned(wire0[(4'h9):(2'h3)]);
            end
          else
            begin
              reg10 <= (wire3 <= (forvar7 ?
                  (~^$unsigned((wire1 ^~ reg13))) : wire3[(3'h5):(2'h2)]));
              reg11 <= reg6[(2'h2):(2'h2)];
              reg14 = $signed($signed(reg11));
              reg15 <= (~&(wire3[(5'h11):(4'h8)] ?
                  wire3 : ({(^~reg12)} ? {(-wire1)} : reg9)));
            end
          if (($unsigned((~{$unsigned(reg5)})) << $signed((+($signed(wire1) ?
              wire3 : (wire2 ? reg15 : reg5))))))
            begin
              reg16 <= reg8[(3'h4):(2'h2)];
            end
          else
            begin
              reg16 <= $signed(reg9);
              reg17 <= $unsigned(wire1);
              reg18 <= (-$unsigned(((-reg9[(1'h0):(1'h0)]) ~^ (^~reg8[(3'h4):(2'h3)]))));
              reg19 <= $signed(reg17[(1'h1):(1'h0)]);
              reg20 = $signed(({($signed(reg10) <<< $unsigned(reg6))} | (~(^~reg17))));
            end
        end
      reg21 <= (~&(!reg14));
    end
  always
    @(posedge clk) begin
      reg22 <= $unsigned((8'hb3));
      reg23 <= (|$signed(reg11[(4'hb):(4'h8)]));
    end
  module24 #() modinst514 (wire513, clk, reg16, reg22, wire1, reg17, reg11);
  module145 #() modinst516 (wire515, clk, wire1, reg11, reg8, wire3);
  module30 #() modinst518 (wire517, clk, reg10, wire1, reg19, reg23, wire513);
  assign wire519 = $signed($signed($unsigned(reg5[(4'ha):(3'h6)])));
  assign wire520 = $unsigned($unsigned((8'hba)));
  module145 #() modinst522 (wire521, clk, reg17, wire513, reg10, reg13);
  always
    @(posedge clk) begin
      reg523 <= (&reg8);
    end
  always
    @(posedge clk) begin
      if ((~&((-$signed((reg21 ? wire3 : wire517))) ?
          (!$signed(wire515)) : $signed($unsigned((wire3 >= wire517))))))
        begin
          reg524 <= $unsigned(reg11[(1'h0):(1'h0)]);
          reg525 <= {(reg13 && ((wire4[(3'h5):(3'h5)] ?
                  $signed(reg13) : (~&reg19)) | reg523)),
              (8'ha6)};
          reg526 <= reg524[(4'he):(4'hd)];
          reg527 <= $unsigned((&(~{(reg19 ? reg524 : wire1)})));
          reg528 <= ((($signed($unsigned(reg5)) ?
                  (~|(reg5 ? reg22 : wire0)) : reg526[(1'h1):(1'h0)]) ?
              (((reg8 ? reg21 : reg13) - (|reg19)) ?
                  reg525 : ($signed((8'hb6)) != ((8'hb2) & wire3))) : {wire515,
                  reg16}) ~^ ($unsigned((-(8'hbd))) ?
              ($unsigned($signed(reg16)) >> (reg22 ?
                  $unsigned(reg527) : (reg5 ?
                      (7'h44) : wire2))) : ($signed((^~reg523)) & {$unsigned(wire520),
                  $unsigned(reg10)})));
        end
      else
        begin
          reg524 <= ({$unsigned((~|(-wire3)))} ?
              $unsigned((&wire515[(1'h1):(1'h1)])) : (reg21 >>> (8'hb3)));
          for (forvar525 = (1'h0); (forvar525 < (2'h2)); forvar525 = (forvar525 + (1'h1)))
            begin
              reg526 <= $signed(wire515[(3'h7):(3'h5)]);
              reg529 = wire515;
            end
          for (forvar530 = (1'h0); (forvar530 < (2'h2)); forvar530 = (forvar530 + (1'h1)))
            begin
              reg531 <= {(wire520[(1'h0):(1'h0)] ?
                      (({reg15, reg21} ?
                          (reg526 == reg12) : reg11[(4'hf):(4'hb)]) - $signed(wire1[(4'h8):(1'h0)])) : reg523)};
              reg532 <= ($signed((8'hac)) << (wire521[(3'h4):(1'h1)] ?
                  ($unsigned((wire4 <= reg526)) ^~ reg525[(1'h0):(1'h0)]) : {reg15[(1'h0):(1'h0)],
                      ((^reg524) ? $signed(reg524) : (~|(8'hac)))}));
              reg533 <= $signed($unsigned({$unsigned($unsigned(wire517))}));
              reg534 = reg527[(4'he):(1'h1)];
              reg535 <= ($unsigned(forvar525[(2'h3):(1'h1)]) >> reg5);
            end
        end
      if ($signed(reg12[(1'h0):(1'h0)]))
        begin
          if ({{($signed((wire520 << wire0)) ? wire1[(4'hd):(1'h1)] : reg6),
                  $signed((reg15[(2'h2):(1'h1)] << $signed(wire0)))},
              ((7'h43) ?
                  (|($unsigned(wire513) >> (reg16 < reg532))) : reg525[(1'h1):(1'h1)])})
            begin
              reg536 <= reg529[(2'h3):(1'h0)];
              reg537 <= ((^(~|reg5)) > reg16[(5'h10):(1'h1)]);
              reg538 <= (~|(-$unsigned(reg17)));
              reg539 <= $unsigned((&(~|(reg529 ~^ {wire513, (8'haa)}))));
              reg540 = $unsigned({(((reg536 ? reg23 : reg526) ?
                          (8'hbf) : reg12[(3'h4):(2'h2)]) ?
                      ($unsigned(reg526) ?
                          $signed(reg19) : $signed(reg5)) : (^reg10)),
                  ({(reg17 ?
                          wire1 : forvar530)} ^~ $unsigned($unsigned(reg539)))});
            end
          else
            begin
              reg540 = {$unsigned(wire519), reg529};
              reg541 <= wire513[(5'h10):(1'h0)];
            end
        end
      else
        begin
          for (forvar536 = (1'h0); (forvar536 < (1'h0)); forvar536 = (forvar536 + (1'h1)))
            begin
              reg540 = $unsigned(reg23);
              reg541 <= forvar536;
              reg542 = (|(!(($signed(reg532) || $unsigned(reg19)) << wire520[(3'h6):(2'h2)])));
            end
          for (forvar543 = (1'h0); (forvar543 < (1'h0)); forvar543 = (forvar543 + (1'h1)))
            begin
              reg544 <= (~^reg534[(1'h1):(1'h0)]);
              reg545 <= (((reg533 | reg536[(3'h4):(1'h0)]) > {$unsigned(reg532[(4'hc):(4'h9)])}) ^~ ((+((^~reg533) ?
                  reg533[(2'h2):(2'h2)] : reg535)) << (reg535[(2'h3):(2'h3)] >> $unsigned($unsigned((8'h9c))))));
              reg546 <= (|((^~$signed((reg21 ?
                  reg532 : (8'hb7)))) <= $signed((-$signed((8'hbe))))));
              reg547 <= (((7'h44) - $unsigned($unsigned(reg537[(2'h2):(1'h0)]))) ?
                  wire3[(4'ha):(3'h4)] : (-(reg546 ?
                      $unsigned(forvar536[(3'h6):(2'h2)]) : ((^~wire517) && (wire521 ?
                          forvar530 : forvar536)))));
              reg548 <= reg23;
            end
        end
      reg549 <= ({$signed(reg13[(4'hb):(3'h4)]),
          forvar543} ^~ (reg525[(1'h1):(1'h1)] << $signed(((reg11 ?
          reg539 : reg21) ~^ (|reg532)))));
      for (forvar550 = (1'h0); (forvar550 < (1'h1)); forvar550 = (forvar550 + (1'h1)))
        begin
          reg551 <= $unsigned($signed($unsigned($signed(((8'hb7) ?
              reg23 : reg524)))));
          reg552 = wire2[(4'ha):(4'ha)];
        end
    end
  always
    @(posedge clk) begin
      reg553 <= reg535[(3'h7):(3'h5)];
      reg554 <= reg6[(3'h4):(3'h4)];
      reg555 <= ((~^((^~(8'hb5)) <= $unsigned($signed(reg554)))) ?
          wire513 : (reg525[(2'h2):(1'h1)] == (-reg525)));
      reg556 <= $signed(((($unsigned(reg5) >= (~(8'ha6))) ?
              $signed(reg547[(3'h6):(3'h6)]) : $signed({wire521})) ?
          ((reg553[(3'h6):(3'h6)] ?
              reg8[(1'h1):(1'h0)] : $unsigned(reg538)) * (!reg537)) : ($signed((reg16 >> (8'ha5))) >> (8'ha8))));
      reg557 <= $unsigned(((~|reg541[(4'ha):(4'h8)]) ?
          $signed($signed(reg545)) : reg555));
    end
  assign wire558 = wire521[(2'h2):(1'h0)];
  module30 #() modinst560 (wire559, clk, reg6, reg8, reg555, reg548, reg22);
  always
    @(posedge clk) begin
      if (reg532[(2'h3):(1'h1)])
        begin
          reg561 = $signed(((~&wire1[(1'h1):(1'h1)]) ~^ $unsigned((reg541 ?
              {reg535} : $signed(reg6)))));
          for (forvar562 = (1'h0); (forvar562 < (2'h3)); forvar562 = (forvar562 + (1'h1)))
            begin
              reg563 <= wire4;
            end
          reg564 <= reg557;
          for (forvar565 = (1'h0); (forvar565 < (3'h4)); forvar565 = (forvar565 + (1'h1)))
            begin
              reg566 <= $unsigned(reg533);
              reg567 <= ($signed($signed($signed($signed(wire513)))) ?
                  $unsigned({$signed($unsigned(reg528)),
                      ((~^wire519) ?
                          $signed(reg524) : ((8'hac) ^~ reg554))}) : $signed(((((8'hac) | reg16) ?
                      (~|wire1) : reg563) ^~ ($signed(wire513) ^ (wire1 ?
                      reg16 : (7'h41))))));
              reg568 = reg564[(3'h5):(2'h3)];
            end
        end
      else
        begin
          reg562 <= $signed(((8'hb2) ? reg8 : (~reg531[(1'h0):(1'h0)])));
          reg563 <= (&$unsigned($unsigned(reg531)));
        end
      reg569 <= ((8'hba) ?
          forvar562 : $signed((reg537[(1'h1):(1'h0)] ?
              reg561 : $unsigned(reg564[(5'h13):(5'h11)]))));
      if ($signed($signed(((reg527 ?
          reg12[(1'h0):(1'h0)] : reg5) ^ ($signed(reg535) ?
          wire2[(2'h3):(2'h2)] : $unsigned(reg536))))))
        begin
          reg570 <= ($unsigned({(8'h9c), (|reg566[(1'h0):(1'h0)])}) ?
              (+({$unsigned((8'hae)),
                  $signed(reg539)} ^ (~&wire4[(4'h8):(3'h6)]))) : (8'ha8));
          if (((wire2 ?
              ((|(reg546 << reg10)) > (~reg567[(1'h0):(1'h0)])) : $signed($unsigned(reg532))) ^ $signed(($unsigned($unsigned(reg19)) * $signed(reg567)))))
            begin
              reg571 <= wire1;
              reg572 <= $unsigned(reg5);
            end
          else
            begin
              reg571 <= wire520[(4'h8):(3'h6)];
              reg572 <= $signed((reg563 * $signed($unsigned((!reg526)))));
            end
        end
      else
        begin
          reg570 <= ((+reg23[(2'h3):(2'h2)]) >> $signed((reg535[(2'h2):(2'h2)] ?
              $signed(((8'ha0) ? wire515 : (8'hb9))) : $signed(reg569))));
          reg571 <= reg555[(4'hf):(3'h7)];
          reg572 <= $signed(($unsigned(reg10) ?
              $unsigned((wire559 ?
                  (reg533 ?
                      reg546 : reg537) : $unsigned(wire558))) : (~&(!reg545[(5'h11):(4'h8)]))));
          for (forvar573 = (1'h0); (forvar573 < (2'h3)); forvar573 = (forvar573 + (1'h1)))
            begin
              reg574 <= ($unsigned({$signed((reg547 > (8'hab)))}) | {$signed(reg537[(2'h2):(2'h2)])});
              reg575 <= wire4;
            end
          for (forvar576 = (1'h0); (forvar576 < (2'h3)); forvar576 = (forvar576 + (1'h1)))
            begin
              reg577 <= $signed((|reg535[(3'h4):(1'h0)]));
            end
        end
      if ({$unsigned($unsigned(reg6[(3'h6):(3'h4)])),
          $signed((~|(reg21[(3'h5):(1'h1)] ?
              $unsigned((8'ha0)) : (reg6 ? reg22 : reg23))))})
        begin
          reg578 <= $signed((~{{$unsigned(wire520)}}));
          reg579 = {reg5[(1'h1):(1'h1)]};
          for (forvar580 = (1'h0); (forvar580 < (1'h0)); forvar580 = (forvar580 + (1'h1)))
            begin
              reg581 <= (~^reg535);
              reg582 <= forvar580;
              reg583 <= $signed(reg574[(4'h9):(2'h2)]);
              reg584 <= reg547[(3'h6):(3'h4)];
            end
        end
      else
        begin
          reg579 = $signed($unsigned(((reg545 ?
                  (reg16 ? reg533 : reg526) : forvar576) ?
              reg549[(3'h7):(1'h1)] : $unsigned(reg8))));
          for (forvar580 = (1'h0); (forvar580 < (1'h1)); forvar580 = (forvar580 + (1'h1)))
            begin
              reg581 <= (&reg581);
              reg582 <= reg528;
              reg583 <= (reg12[(2'h2):(2'h2)] ? wire0 : $signed((8'ha3)));
            end
          reg584 <= reg568[(4'h9):(2'h2)];
        end
      reg585 <= reg566[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg586 <= (((~^reg569) ?
              $signed((-$unsigned(reg564))) : (reg531 ?
                  $signed((8'hbb)) : ($signed(reg19) ?
                      (wire519 ? reg531 : wire521) : (reg528 ?
                          reg574 : reg574)))) ?
          ((-$unsigned((reg525 >= reg22))) ?
              (reg571 > ((reg575 < reg535) - $unsigned(reg524))) : reg8) : (|$signed((~&(!reg569)))));
    end
  always
    @(posedge clk) begin
      reg587 <= (8'hab);
      for (forvar588 = (1'h0); (forvar588 < (3'h4)); forvar588 = (forvar588 + (1'h1)))
        begin
          reg589 = (!$unsigned($unsigned(((^~reg21) ?
              (+reg547) : reg563[(3'h5):(1'h1)]))));
          reg590 <= reg557;
          reg591 <= (({(+(reg571 ? reg544 : reg532))} ?
              $signed(reg583) : $signed(reg584[(4'h8):(3'h5)])) || (~|reg590));
          reg592 <= {{$unsigned(reg563), $signed($unsigned((!reg556)))},
              ((~^reg533) >> ((reg12 ? reg541 : (-(8'h9d))) ?
                  $unsigned(reg537[(1'h0):(1'h0)]) : ((reg577 ?
                      reg21 : reg569) && wire1)))};
          reg593 <= $unsigned(reg549);
        end
      for (forvar594 = (1'h0); (forvar594 < (1'h0)); forvar594 = (forvar594 + (1'h1)))
        begin
          reg595 <= $unsigned((reg22 == ((reg537 - reg19[(3'h4):(1'h1)]) || reg549[(3'h4):(1'h1)])));
          if (reg532[(2'h2):(1'h1)])
            begin
              reg596 <= (|(reg11[(1'h0):(1'h0)] | ($unsigned((reg8 ?
                  reg15 : wire519)) == (-(reg545 ? (8'haf) : reg581)))));
              reg597 <= $unsigned(((reg531[(3'h5):(1'h0)] ?
                      ($unsigned(reg532) ?
                          $signed(reg562) : $unsigned(reg546)) : reg526[(3'h7):(2'h3)]) ?
                  wire521 : reg564[(1'h0):(1'h0)]));
              reg598 <= (~&reg527);
            end
          else
            begin
              reg596 <= (|(~{$unsigned((reg548 ? reg566 : reg587))}));
            end
          if ($unsigned((^$unsigned(($signed((8'hb2)) ?
              (+wire4) : $unsigned(reg598))))))
            begin
              reg599 <= reg18;
              reg600 = reg12;
              reg601 <= $signed((|reg547));
              reg602 <= (^~(($unsigned($unsigned(wire0)) ?
                  $signed($unsigned(reg571)) : $unsigned((^reg582))) * ((reg12[(1'h0):(1'h0)] ?
                      $signed(wire520) : reg557[(2'h3):(2'h2)]) ?
                  wire3[(1'h1):(1'h1)] : $unsigned($unsigned(reg13)))));
            end
          else
            begin
              reg599 <= $signed((-($signed(((8'ha5) ~^ (8'hbc))) >> (~&(wire3 ?
                  reg587 : reg11)))));
              reg601 <= reg582;
              reg603 = wire2;
            end
          reg604 <= reg551[(3'h7):(1'h1)];
        end
      reg605 <= reg575;
      reg606 <= (-reg17);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module24  (y, clk, wire25, wire26, wire27, wire28, wire29);
  output wire [(32'h239):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire25;
  input wire [(4'h8):(1'h0)] wire26;
  input wire [(4'hb):(1'h0)] wire27;
  input wire [(5'h14):(1'h0)] wire28;
  input wire signed [(5'h12):(1'h0)] wire29;
  wire [(5'h13):(1'h0)] wire479;
  wire signed [(5'h14):(1'h0)] wire414;
  wire signed [(3'h6):(1'h0)] wire387;
  wire [(4'hc):(1'h0)] wire290;
  wire [(5'h14):(1'h0)] wire143;
  wire [(5'h13):(1'h0)] wire471;
  wire [(5'h10):(1'h0)] wire473;
  wire signed [(3'h5):(1'h0)] wire474;
  wire signed [(5'h11):(1'h0)] wire475;
  wire signed [(4'h9):(1'h0)] wire476;
  wire signed [(5'h11):(1'h0)] wire477;
  wire [(5'h11):(1'h0)] wire481;
  wire [(5'h11):(1'h0)] wire482;
  wire [(3'h7):(1'h0)] wire484;
  reg signed [(4'hc):(1'h0)] reg512 = (1'h0);
  reg [(4'h9):(1'h0)] reg511 = (1'h0);
  reg [(3'h4):(1'h0)] reg510 = (1'h0);
  reg [(4'hc):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg506 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg505 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg504 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg503 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg502 = (1'h0);
  reg [(4'hb):(1'h0)] reg500 = (1'h0);
  reg [(5'h10):(1'h0)] reg498 = (1'h0);
  reg [(2'h3):(1'h0)] reg497 = (1'h0);
  reg [(2'h3):(1'h0)] reg495 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg494 = (1'h0);
  reg [(5'h10):(1'h0)] reg493 = (1'h0);
  reg [(3'h4):(1'h0)] reg492 = (1'h0);
  reg [(5'h14):(1'h0)] reg491 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg486 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg417 = (1'h0);
  reg [(4'hf):(1'h0)] reg416 = (1'h0);
  reg [(3'h6):(1'h0)] reg293 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg389 = (1'h0);
  reg [(4'h8):(1'h0)] reg508 = (1'h0);
  reg [(4'hb):(1'h0)] reg507 = (1'h0);
  reg [(4'hd):(1'h0)] forvar501 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg499 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg496 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg490 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg489 = (1'h0);
  reg [(4'hf):(1'h0)] reg488 = (1'h0);
  reg [(5'h11):(1'h0)] forvar487 = (1'h0);
  reg signed [(4'he):(1'h0)] reg292 = (1'h0);
  assign y = {wire479,
                 wire414,
                 wire387,
                 wire290,
                 wire143,
                 wire471,
                 wire473,
                 wire474,
                 wire475,
                 wire476,
                 wire477,
                 wire481,
                 wire482,
                 wire484,
                 reg512,
                 reg511,
                 reg510,
                 reg509,
                 reg506,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 reg500,
                 reg498,
                 reg497,
                 reg495,
                 reg494,
                 reg493,
                 reg492,
                 reg491,
                 reg486,
                 reg417,
                 reg416,
                 reg293,
                 reg389,
                 reg508,
                 reg507,
                 forvar501,
                 reg499,
                 reg496,
                 reg490,
                 reg489,
                 reg488,
                 forvar487,
                 reg292,
                 (1'h0)};
  module30 #() modinst144 (wire143, clk, wire25, wire29, wire27, wire26, wire28);
  module145 #() modinst291 (.clk(clk), .wire149(wire27), .wire146(wire29), .y(wire290), .wire147(wire25), .wire148(wire28));
  always
    @(posedge clk) begin
      reg292 = $signed(wire290[(1'h0):(1'h0)]);
      reg293 <= reg292[(2'h2):(1'h0)];
    end
  module294 #() modinst388 (.wire296(wire29), .wire298(wire143), .wire297(wire27), .wire295(wire290), .clk(clk), .y(wire387));
  always
    @(posedge clk) begin
      reg389 <= $unsigned((^~reg293[(1'h1):(1'h0)]));
    end
  module390 #() modinst415 (.wire391(wire27), .wire393(wire25), .y(wire414), .wire394(reg389), .clk(clk), .wire392(wire290));
  always
    @(posedge clk) begin
      reg416 <= ((^(wire414[(1'h0):(1'h0)] != ({wire29} <= reg293))) > wire25[(4'hf):(1'h0)]);
      reg417 <= wire29;
    end
  module418 #() modinst472 (wire471, clk, reg293, wire27, wire414, wire29, wire290);
  assign wire473 = (wire27[(1'h0):(1'h0)] ?
                       $unsigned((((~&wire27) && (reg417 ? wire26 : reg416)) ?
                           $signed((-wire26)) : $unsigned(wire26[(3'h6):(1'h1)]))) : (8'hb5));
  assign wire474 = $signed($signed((!($unsigned(wire27) ?
                       wire29 : (wire473 >> reg293)))));
  assign wire475 = wire26;
  assign wire476 = (wire290 == (wire25[(5'h13):(5'h12)] > $signed(($unsigned(wire29) ?
                       $signed(wire474) : (&wire26)))));
  module390 #() modinst478 (.wire393(reg417), .y(wire477), .wire392(wire143), .wire394(wire25), .clk(clk), .wire391(wire414));
  module418 #() modinst480 (wire479, clk, wire414, wire476, wire29, wire25, wire290);
  assign wire481 = (~^(wire476 ? $signed(wire26) : {wire473}));
  module30 #() modinst483 (.wire33(wire28), .wire32(wire25), .wire31(wire414), .clk(clk), .y(wire482), .wire35(wire143), .wire34(reg416));
  module390 #() modinst485 (.wire394(wire25), .clk(clk), .wire393(wire473), .wire391(reg389), .y(wire484), .wire392(wire28));
  always
    @(posedge clk) begin
      reg486 <= (8'hbc);
      for (forvar487 = (1'h0); (forvar487 < (3'h4)); forvar487 = (forvar487 + (1'h1)))
        begin
          reg488 = $unsigned(wire25);
          if ((wire481 & $signed(($unsigned($signed(wire477)) ?
              wire471 : $unsigned(wire479[(5'h10):(4'hb)])))))
            begin
              reg489 = wire471[(4'h9):(1'h0)];
              reg490 = ((reg486[(3'h6):(3'h5)] ?
                      $signed(reg488) : wire479[(3'h6):(1'h1)]) ?
                  {((~|((8'ha7) ? wire479 : wire290)) ?
                          $unsigned($signed(wire290)) : wire481[(2'h3):(2'h2)])} : ((~&{((8'h9c) ?
                              wire28 : wire143)}) ?
                      $unsigned($unsigned((^~wire473))) : $signed((((8'hbc) ?
                          wire473 : reg416) || wire29))));
            end
          else
            begin
              reg491 <= $unsigned(((8'hbb) ?
                  ((~&$signed(wire471)) ?
                      $unsigned(wire477[(4'he):(4'ha)]) : (&(-wire473))) : {((wire482 ?
                              wire482 : (8'ha6)) ?
                          wire481[(4'h9):(2'h2)] : {(8'hb1), wire26})}));
            end
          reg492 <= (-$unsigned((wire471 | (reg416 >> (wire477 >> wire477)))));
          reg493 <= (~{$signed(reg492[(2'h3):(1'h0)]),
              $unsigned(({wire471} <<< $signed(wire482)))});
        end
      if ((wire477[(2'h2):(1'h0)] ?
          ($signed($unsigned((~^reg488))) ?
              reg416 : wire28) : wire481[(4'h9):(3'h5)]))
        begin
          reg494 <= reg293[(1'h0):(1'h0)];
          reg495 <= ($signed(wire25) | (wire29 ?
              ($signed(reg493[(4'h8):(2'h2)]) < {wire484[(1'h0):(1'h0)]}) : $signed((wire482 >>> (~wire29)))));
          reg496 = $signed($unsigned((~|$unsigned(reg416[(2'h2):(2'h2)]))));
          reg497 <= (wire484 ? (&{$unsigned({reg491, reg417})}) : reg490);
          reg498 <= $unsigned({(-($unsigned((8'h9d)) ?
                  (wire29 ? wire482 : wire476) : (^~wire482))),
              $signed(wire414[(5'h12):(3'h6)])});
        end
      else
        begin
          reg494 <= wire28;
          reg495 <= wire290;
          reg496 = ($unsigned($signed((!reg497))) ^ (^$unsigned(reg498[(4'hb):(3'h6)])));
          reg497 <= wire484;
        end
      reg499 = (~|($signed(reg493) != (~^wire476[(1'h0):(1'h0)])));
    end
  always
    @(posedge clk) begin
      reg500 <= (~&(8'hbe));
      for (forvar501 = (1'h0); (forvar501 < (2'h2)); forvar501 = (forvar501 + (1'h1)))
        begin
          if (($unsigned(($signed({forvar501, wire25}) | {{wire414,
                  wire143}})) <<< {((8'hb9) + wire29[(4'hb):(3'h6)]), wire479}))
            begin
              reg502 <= forvar501[(3'h4):(2'h3)];
              reg503 <= (((~&((^~(8'hab)) <= $signed((7'h42)))) & ({$signed(wire476)} ?
                      $signed((^wire471)) : (|(&reg416)))) ?
                  $signed(wire474) : ({(reg495[(2'h3):(2'h2)] ?
                              $unsigned(wire143) : ((8'hb4) >> wire477))} ?
                      {$signed(reg498[(3'h7):(1'h0)]),
                          (((7'h40) || wire474) ~^ reg417[(1'h1):(1'h0)])} : ($signed($signed((8'haf))) < ((+reg416) ?
                          (!wire28) : $signed(reg493)))));
              reg504 <= $unsigned(wire475[(2'h2):(2'h2)]);
              reg505 <= (+$signed($unsigned($unsigned($signed((8'ha3))))));
              reg506 <= $unsigned(wire476);
            end
          else
            begin
              reg502 <= $signed($signed({(reg502[(3'h4):(1'h1)] - $signed(reg491)),
                  $signed(reg503)}));
              reg503 <= ({reg502[(3'h4):(2'h3)],
                      $signed($signed($signed((8'ha6))))} ?
                  ((8'hbe) | wire290) : $unsigned($unsigned($unsigned((reg495 ?
                      wire475 : reg417)))));
              reg504 <= reg497[(1'h0):(1'h0)];
              reg505 <= reg497;
              reg506 <= $unsigned(wire481);
            end
        end
      if (reg505)
        begin
          reg507 = $unsigned(({$signed((~wire482)), reg293} & reg502));
          reg508 = ($signed($unsigned($unsigned((wire477 != reg505)))) == ($unsigned((^(reg417 >> wire387))) ?
              $signed(((~&wire482) ? $signed(reg495) : reg503)) : ((reg494 ?
                      (wire479 >= reg503) : (wire481 ? wire27 : wire28)) ?
                  (wire471 ? (!wire29) : reg491[(2'h2):(1'h1)]) : ((reg495 ?
                          reg493 : reg506) ?
                      (reg500 ^ wire473) : (reg494 ? reg500 : reg500)))));
          reg509 <= ($signed($unsigned(($signed(reg389) ?
              $signed(wire414) : {reg504,
                  wire387}))) != (reg493[(1'h0):(1'h0)] & ($unsigned((reg493 >= wire477)) ?
              (+forvar501) : forvar501[(2'h3):(2'h2)])));
        end
      else
        begin
          if (wire475)
            begin
              reg509 <= (reg498[(4'h8):(3'h6)] ?
                  (!$signed(reg498[(4'hd):(3'h7)])) : wire471);
              reg510 <= (wire476 ^ ($signed($signed((!reg505))) ?
                  (8'hb1) : (reg495[(1'h0):(1'h0)] && wire482[(5'h11):(1'h0)])));
              reg511 <= forvar501[(1'h0):(1'h0)];
            end
          else
            begin
              reg509 <= $unsigned((reg492[(2'h3):(1'h1)] >> ($unsigned((reg510 ?
                  wire475 : wire414)) || (~^{wire28, wire290}))));
            end
          reg512 <= $unsigned($signed(reg506));
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module418
#(parameter param469 = {((&(8'hbe)) ? ((^(~^(8'ha4))) >> ((~^(8'ha2)) ^ ((8'hac) ? (8'ha2) : (8'haf)))) : ({(7'h42)} < ({(8'h9d)} & (8'hb5)))), (!(-(-((8'ha6) ? (8'hab) : (7'h42)))))}, 
parameter param470 = {(8'hb8)})
(y, clk, wire423, wire422, wire421, wire420, wire419);
  output wire [(32'h1f0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h6):(1'h0)] wire423;
  input wire [(4'h9):(1'h0)] wire422;
  input wire [(3'h6):(1'h0)] wire421;
  input wire [(4'ha):(1'h0)] wire420;
  input wire [(4'h9):(1'h0)] wire419;
  wire signed [(3'h5):(1'h0)] wire468;
  wire [(2'h2):(1'h0)] wire453;
  reg signed [(3'h5):(1'h0)] reg467 = (1'h0);
  reg [(5'h14):(1'h0)] reg466 = (1'h0);
  reg [(5'h11):(1'h0)] reg465 = (1'h0);
  reg [(5'h12):(1'h0)] reg464 = (1'h0);
  reg [(5'h10):(1'h0)] reg463 = (1'h0);
  reg [(3'h7):(1'h0)] reg462 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg461 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg460 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg459 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg455 = (1'h0);
  reg signed [(4'he):(1'h0)] reg454 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg452 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg451 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg450 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg449 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg448 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg447 = (1'h0);
  reg [(4'ha):(1'h0)] reg445 = (1'h0);
  reg [(4'hc):(1'h0)] reg444 = (1'h0);
  reg [(4'hc):(1'h0)] reg443 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg442 = (1'h0);
  reg [(3'h7):(1'h0)] reg441 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg440 = (1'h0);
  reg [(2'h3):(1'h0)] reg437 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg436 = (1'h0);
  reg [(4'ha):(1'h0)] reg435 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg434 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg433 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg432 = (1'h0);
  reg [(3'h4):(1'h0)] reg431 = (1'h0);
  reg [(3'h7):(1'h0)] reg430 = (1'h0);
  reg [(5'h10):(1'h0)] reg427 = (1'h0);
  reg [(2'h2):(1'h0)] reg425 = (1'h0);
  reg [(3'h5):(1'h0)] reg458 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar457 = (1'h0);
  reg [(2'h3):(1'h0)] forvar456 = (1'h0);
  reg [(5'h10):(1'h0)] reg446 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar439 = (1'h0);
  reg [(4'h9):(1'h0)] forvar438 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar429 = (1'h0);
  reg [(4'hf):(1'h0)] reg428 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg426 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar424 = (1'h0);
  assign y = {wire468,
                 wire453,
                 reg467,
                 reg466,
                 reg465,
                 reg464,
                 reg463,
                 reg462,
                 reg461,
                 reg460,
                 reg459,
                 reg455,
                 reg454,
                 reg452,
                 reg451,
                 reg450,
                 reg449,
                 reg448,
                 reg447,
                 reg445,
                 reg444,
                 reg443,
                 reg442,
                 reg441,
                 reg440,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg433,
                 reg432,
                 reg431,
                 reg430,
                 reg427,
                 reg425,
                 reg458,
                 forvar457,
                 forvar456,
                 reg446,
                 forvar439,
                 forvar438,
                 forvar429,
                 reg428,
                 reg426,
                 forvar424,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar424 = (1'h0); (forvar424 < (1'h1)); forvar424 = (forvar424 + (1'h1)))
        begin
          reg425 <= (($unsigned(($unsigned(wire420) ?
                  (forvar424 + wire423) : $unsigned(forvar424))) <<< (((forvar424 ?
                  wire421 : wire419) ~^ wire420) * $signed((^~wire419)))) ?
              (|(&$signed(wire421[(2'h2):(1'h1)]))) : ((wire419[(2'h3):(1'h0)] + $unsigned((wire423 | wire420))) != $signed(($unsigned(wire419) & $unsigned(wire422)))));
          reg426 = $signed(((~(forvar424 + $unsigned(wire419))) & (+((wire421 ?
              wire422 : (8'ha3)) && (wire421 ? (8'hb1) : reg425)))));
          reg427 <= (8'hb2);
          reg428 = (reg426[(3'h7):(2'h2)] ?
              ($unsigned(((wire422 ?
                  reg425 : reg426) && wire420[(4'ha):(4'ha)])) + (wire419[(1'h0):(1'h0)] ?
                  forvar424[(4'h8):(2'h2)] : wire420[(1'h0):(1'h0)])) : $unsigned(((~&(!forvar424)) == (reg425 == (~^(8'hab))))));
          for (forvar429 = (1'h0); (forvar429 < (2'h2)); forvar429 = (forvar429 + (1'h1)))
            begin
              reg430 <= reg427[(3'h4):(2'h2)];
            end
        end
      reg431 <= $unsigned($unsigned(({$signed(reg426), reg430} ?
          wire419 : $signed(wire421[(1'h0):(1'h0)]))));
      reg432 <= reg428;
      reg433 <= (~((~^(forvar429[(3'h6):(3'h4)] ?
          (^~(8'haf)) : $unsigned(wire421))) << forvar429));
    end
  always
    @(posedge clk) begin
      reg434 <= $unsigned((($unsigned($signed(wire420)) ?
              ({reg432, (8'h9c)} ?
                  (~wire419) : $signed(reg431)) : $unsigned((reg427 >= wire423))) ?
          $unsigned((reg430[(3'h5):(1'h1)] ?
              $signed((8'hbe)) : reg430[(3'h7):(1'h1)])) : (^$signed((~^(7'h40))))));
      reg435 <= ((wire421 ? {$unsigned(reg431)} : $unsigned(wire422)) ?
          $signed($signed((reg427 ?
              (wire423 ?
                  (8'haf) : wire422) : (reg425 <<< wire422)))) : reg432[(4'ha):(4'h9)]);
      reg436 <= $signed($signed(wire423[(1'h1):(1'h0)]));
      reg437 <= reg430;
    end
  always
    @(posedge clk) begin
      for (forvar438 = (1'h0); (forvar438 < (1'h0)); forvar438 = (forvar438 + (1'h1)))
        begin
          for (forvar439 = (1'h0); (forvar439 < (2'h3)); forvar439 = (forvar439 + (1'h1)))
            begin
              reg440 <= (^$unsigned(reg433[(1'h1):(1'h0)]));
              reg441 <= $unsigned($unsigned({(~&(~&(8'ha2))),
                  $unsigned(reg427)}));
              reg442 <= {wire422};
              reg443 <= reg432[(3'h4):(1'h1)];
              reg444 <= $signed(($unsigned(wire420) < $signed($unsigned(reg441[(2'h3):(2'h3)]))));
            end
          if (reg434)
            begin
              reg445 <= (~^({$unsigned((!reg435))} && ($signed((reg425 ?
                      forvar439 : (8'hbf))) ?
                  (8'hbe) : reg436[(3'h5):(2'h2)])));
              reg446 = {$unsigned({$unsigned($signed(reg431))})};
              reg447 <= wire423[(3'h4):(2'h2)];
              reg448 <= {$signed($signed((reg432[(4'hf):(2'h2)] ?
                      (8'ha8) : $signed(reg437)))),
                  (+$signed($unsigned({reg437, (7'h40)})))};
              reg449 <= ($signed(reg431[(1'h0):(1'h0)]) ?
                  $signed(($signed({(8'hb9), reg448}) ?
                      (reg431 ?
                          (~&reg431) : $signed(reg445)) : $signed(reg443[(2'h2):(1'h0)]))) : $signed($unsigned({reg427[(4'h9):(3'h4)],
                      reg443[(3'h5):(1'h1)]})));
            end
          else
            begin
              reg445 <= $unsigned(reg447[(3'h4):(1'h0)]);
              reg447 <= $unsigned(($unsigned($unsigned((reg435 ?
                  reg436 : reg427))) ~^ (wire423 ?
                  reg432[(5'h11):(5'h11)] : (^(reg443 ? wire421 : reg448)))));
            end
          reg450 <= reg441[(2'h2):(1'h0)];
          reg451 <= (~^$unsigned(reg437[(2'h3):(2'h3)]));
          reg452 <= reg449[(2'h2):(2'h2)];
        end
    end
  assign wire453 = $signed(((reg427 ^~ (~&$unsigned((8'h9e)))) ?
                       reg427[(4'hd):(1'h0)] : (((-(8'ha7)) ?
                               reg448 : $unsigned(reg437)) ?
                           $unsigned($unsigned(reg432)) : (reg434 >= $signed((8'ha9))))));
  always
    @(posedge clk) begin
      reg454 <= $signed(((|$signed(reg445)) & (8'hbd)));
      reg455 <= {(~&$signed(($unsigned(reg454) ?
              $unsigned(reg431) : ((8'hae) & (8'hac)))))};
      for (forvar456 = (1'h0); (forvar456 < (1'h1)); forvar456 = (forvar456 + (1'h1)))
        begin
          for (forvar457 = (1'h0); (forvar457 < (2'h3)); forvar457 = (forvar457 + (1'h1)))
            begin
              reg458 = reg447[(1'h0):(1'h0)];
              reg459 <= {(($unsigned(reg449) >= ({(8'ha3),
                          reg449} == (&reg451))) ?
                      ($unsigned(((8'h9e) & wire422)) <<< (wire420[(3'h4):(1'h1)] ?
                          $unsigned(reg450) : ((8'ha6) >= (8'ha8)))) : (-reg448))};
              reg460 <= $signed($unsigned((({(8'ha7), reg442} ?
                      (8'ha9) : $unsigned(reg443)) ?
                  (~&(wire423 * forvar456)) : reg431)));
            end
          reg461 <= ({$unsigned(reg449)} < wire421);
          if ($unsigned(((~&wire423) < {(reg461[(2'h3):(1'h1)] - (reg444 ?
                  reg461 : reg448))})))
            begin
              reg462 <= {$unsigned(((reg436 ?
                          (reg432 ? forvar456 : reg454) : reg432) ?
                      wire422 : ((7'h43) <<< wire423[(3'h4):(2'h2)]))),
                  $unsigned($unsigned((^$signed(reg425))))};
              reg463 <= (~&(~$signed((reg441 >= ((8'ha3) ?
                  reg441 : wire420)))));
              reg464 <= (8'ha4);
              reg465 <= $signed(reg436);
            end
          else
            begin
              reg462 <= reg460[(4'h8):(3'h4)];
              reg463 <= {reg425[(2'h2):(1'h0)], reg430};
            end
          reg466 <= (~^(-{(+(reg440 ^ reg462)),
              $signed(((7'h41) ? reg431 : reg454))}));
          reg467 <= reg451;
        end
    end
  assign wire468 = ($signed(reg449[(1'h1):(1'h1)]) * reg432[(1'h1):(1'h0)]);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module390  (y, clk, wire394, wire393, wire392, wire391);
  output wire [(32'hb8):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h12):(1'h0)] wire394;
  input wire signed [(3'h7):(1'h0)] wire393;
  input wire [(2'h3):(1'h0)] wire392;
  input wire signed [(3'h7):(1'h0)] wire391;
  wire [(5'h10):(1'h0)] wire413;
  wire signed [(5'h15):(1'h0)] wire407;
  wire [(3'h7):(1'h0)] wire406;
  wire [(3'h5):(1'h0)] wire405;
  wire signed [(5'h14):(1'h0)] wire404;
  wire [(4'hc):(1'h0)] wire403;
  reg [(3'h4):(1'h0)] reg412 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg411 = (1'h0);
  reg [(4'hc):(1'h0)] reg410 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg409 = (1'h0);
  reg [(3'h6):(1'h0)] reg402 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg401 = (1'h0);
  reg [(4'hd):(1'h0)] reg400 = (1'h0);
  reg [(5'h13):(1'h0)] reg399 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg397 = (1'h0);
  reg [(4'ha):(1'h0)] reg396 = (1'h0);
  reg [(3'h4):(1'h0)] reg395 = (1'h0);
  reg [(3'h5):(1'h0)] forvar408 = (1'h0);
  reg [(4'h8):(1'h0)] forvar398 = (1'h0);
  assign y = {wire413,
                 wire407,
                 wire406,
                 wire405,
                 wire404,
                 wire403,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg402,
                 reg401,
                 reg400,
                 reg399,
                 reg397,
                 reg396,
                 reg395,
                 forvar408,
                 forvar398,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg395 <= wire393[(3'h7):(3'h7)];
    end
  always
    @(posedge clk) begin
      reg396 <= wire391[(1'h0):(1'h0)];
      reg397 <= ((7'h41) ^~ $signed((~^($signed(reg396) ?
          (reg396 - reg396) : $signed(wire394)))));
    end
  always
    @(posedge clk) begin
      for (forvar398 = (1'h0); (forvar398 < (2'h2)); forvar398 = (forvar398 + (1'h1)))
        begin
          reg399 <= (~$unsigned((~&wire394[(4'hf):(4'hf)])));
        end
    end
  always
    @(posedge clk) begin
      reg400 <= wire392[(2'h3):(2'h3)];
      reg401 <= $unsigned({$signed(reg395[(1'h1):(1'h0)]), reg397});
    end
  always
    @(posedge clk) begin
      reg402 <= (+reg397);
    end
  assign wire403 = wire393;
  assign wire404 = (|(wire394 ? (+{(8'h9f), wire392}) : reg400));
  assign wire405 = ((!$unsigned({$unsigned(reg401)})) ?
                       ({reg400, reg396} ?
                           (|wire404) : (wire391 ?
                               wire403[(4'ha):(3'h6)] : $signed((wire394 ?
                                   reg399 : reg396)))) : $signed(wire403));
  assign wire406 = (wire392[(2'h3):(1'h1)] * wire404[(3'h5):(1'h1)]);
  assign wire407 = {(reg402[(2'h3):(2'h3)] ?
                           ((~&{(8'ha3)}) >= $signed((reg401 ?
                               (7'h42) : wire392))) : reg396),
                       $unsigned({(8'hbd),
                           (reg399 ? ((7'h40) ? reg397 : wire393) : wire391)})};
  always
    @(posedge clk) begin
      for (forvar408 = (1'h0); (forvar408 < (3'h4)); forvar408 = (forvar408 + (1'h1)))
        begin
          reg409 <= (-(!{wire391[(3'h5):(3'h4)]}));
          reg410 <= {wire404,
              $unsigned(((wire407 ^~ (wire393 != reg401)) || {(reg399 ?
                      reg399 : wire393)}))};
        end
      reg411 <= (forvar408[(1'h1):(1'h0)] ?
          (&reg409) : $unsigned(reg410[(2'h3):(2'h2)]));
      reg412 <= ((8'hba) ?
          (((-(reg410 >= wire407)) != reg402[(3'h4):(2'h3)]) ?
              reg395[(2'h3):(1'h0)] : wire405[(3'h4):(1'h1)]) : (~&$unsigned(({reg409} ?
              {reg396} : (reg397 >= reg411)))));
    end
  assign wire413 = (8'hb6);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module294
#(parameter param386 = (&(~^({(-(7'h41)), ((8'ha5) ? (8'hb8) : (8'hbf))} ? (&(!(8'hbe))) : (((8'ha9) ? (8'hbc) : (8'hb2)) ? {(8'ha1), (8'ha0)} : ((8'hb9) ? (8'hb5) : (8'ha9)))))))
(y, clk, wire298, wire297, wire296, wire295);
  output wire [(32'h3f5):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(2'h2):(1'h0)] wire298;
  input wire signed [(4'hb):(1'h0)] wire297;
  input wire signed [(5'h12):(1'h0)] wire296;
  input wire [(4'hc):(1'h0)] wire295;
  wire signed [(3'h5):(1'h0)] wire385;
  wire signed [(2'h2):(1'h0)] wire360;
  wire [(2'h3):(1'h0)] wire338;
  wire [(4'hc):(1'h0)] wire337;
  wire signed [(4'hc):(1'h0)] wire336;
  wire [(4'he):(1'h0)] wire325;
  reg signed [(3'h4):(1'h0)] reg384 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg383 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg382 = (1'h0);
  reg [(3'h4):(1'h0)] reg381 = (1'h0);
  reg [(4'hc):(1'h0)] reg379 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg378 = (1'h0);
  reg [(4'ha):(1'h0)] reg377 = (1'h0);
  reg [(4'hd):(1'h0)] reg376 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg375 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg374 = (1'h0);
  reg [(4'h9):(1'h0)] reg373 = (1'h0);
  reg [(3'h5):(1'h0)] reg372 = (1'h0);
  reg [(5'h11):(1'h0)] reg371 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg369 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg368 = (1'h0);
  reg [(4'hd):(1'h0)] reg367 = (1'h0);
  reg signed [(4'he):(1'h0)] reg365 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg363 = (1'h0);
  reg [(4'ha):(1'h0)] reg362 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg359 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg358 = (1'h0);
  reg [(3'h5):(1'h0)] reg357 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg356 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg355 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg354 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg353 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg351 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg350 = (1'h0);
  reg [(3'h4):(1'h0)] reg344 = (1'h0);
  reg [(5'h15):(1'h0)] reg349 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg348 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg347 = (1'h0);
  reg [(5'h14):(1'h0)] reg346 = (1'h0);
  reg [(4'h8):(1'h0)] reg345 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg343 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg342 = (1'h0);
  reg [(2'h2):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg340 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg339 = (1'h0);
  reg [(3'h7):(1'h0)] reg335 = (1'h0);
  reg [(5'h15):(1'h0)] reg334 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg332 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg331 = (1'h0);
  reg [(3'h6):(1'h0)] reg330 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg328 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg327 = (1'h0);
  reg [(3'h5):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg323 = (1'h0);
  reg [(3'h6):(1'h0)] reg322 = (1'h0);
  reg [(5'h15):(1'h0)] reg319 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg317 = (1'h0);
  reg [(2'h2):(1'h0)] reg315 = (1'h0);
  reg [(4'hd):(1'h0)] reg314 = (1'h0);
  reg [(5'h15):(1'h0)] reg313 = (1'h0);
  reg [(4'h8):(1'h0)] reg312 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg311 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg307 = (1'h0);
  reg [(4'hb):(1'h0)] reg306 = (1'h0);
  reg [(4'hc):(1'h0)] reg305 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg304 = (1'h0);
  reg [(4'hf):(1'h0)] reg303 = (1'h0);
  reg [(4'hd):(1'h0)] reg302 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg301 = (1'h0);
  reg [(2'h2):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg299 = (1'h0);
  reg [(2'h2):(1'h0)] forvar380 = (1'h0);
  reg [(3'h7):(1'h0)] reg370 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg366 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg364 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar361 = (1'h0);
  reg [(4'h8):(1'h0)] forvar352 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar344 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg333 = (1'h0);
  reg [(5'h15):(1'h0)] reg329 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar326 = (1'h0);
  reg [(5'h14):(1'h0)] forvar321 = (1'h0);
  reg [(3'h7):(1'h0)] reg320 = (1'h0);
  reg [(4'he):(1'h0)] reg318 = (1'h0);
  reg [(3'h6):(1'h0)] forvar316 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar310 = (1'h0);
  reg [(5'h11):(1'h0)] reg309 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar301 = (1'h0);
  assign y = {wire385,
                 wire360,
                 wire338,
                 wire337,
                 wire336,
                 wire325,
                 reg384,
                 reg383,
                 reg382,
                 reg381,
                 reg379,
                 reg378,
                 reg377,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg369,
                 reg368,
                 reg367,
                 reg365,
                 reg363,
                 reg362,
                 reg359,
                 reg358,
                 reg357,
                 reg356,
                 reg355,
                 reg354,
                 reg353,
                 reg351,
                 reg350,
                 reg344,
                 reg349,
                 reg348,
                 reg347,
                 reg346,
                 reg345,
                 reg343,
                 reg342,
                 reg341,
                 reg340,
                 reg339,
                 reg335,
                 reg334,
                 reg332,
                 reg331,
                 reg330,
                 reg328,
                 reg327,
                 reg324,
                 reg323,
                 reg322,
                 reg319,
                 reg317,
                 reg315,
                 reg314,
                 reg313,
                 reg312,
                 reg311,
                 reg308,
                 reg307,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg302,
                 reg301,
                 reg300,
                 reg299,
                 forvar380,
                 reg370,
                 reg366,
                 reg364,
                 forvar361,
                 forvar352,
                 forvar344,
                 reg333,
                 reg329,
                 forvar326,
                 forvar321,
                 reg320,
                 reg318,
                 forvar316,
                 forvar310,
                 reg309,
                 forvar301,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg299 <= (-$unsigned(wire297[(1'h0):(1'h0)]));
      reg300 <= (!{wire296});
      if ($signed(reg300[(2'h2):(1'h0)]))
        begin
          reg301 <= {wire295[(2'h2):(2'h2)], wire298[(2'h2):(2'h2)]};
        end
      else
        begin
          for (forvar301 = (1'h0); (forvar301 < (3'h4)); forvar301 = (forvar301 + (1'h1)))
            begin
              reg302 <= (^wire296[(2'h2):(1'h0)]);
              reg303 <= (~({$unsigned(wire295[(4'hb):(4'h9)])} || (+$signed({forvar301}))));
              reg304 <= reg299[(3'h7):(2'h2)];
              reg305 <= wire296;
              reg306 <= reg301;
            end
          if ($unsigned(reg306[(1'h0):(1'h0)]))
            begin
              reg307 <= ((|{{reg306[(1'h0):(1'h0)]}, (^~(^~wire297))}) ?
                  reg301 : ((^(reg302[(3'h5):(3'h4)] ?
                          reg300 : $signed((8'ha5)))) ?
                      (+reg305) : reg301[(4'h9):(1'h0)]));
              reg308 <= $unsigned({(((|(8'hb6)) == forvar301) <<< {$unsigned((8'ha9))}),
                  (^reg300[(2'h2):(1'h0)])});
            end
          else
            begin
              reg309 = forvar301[(1'h0):(1'h0)];
            end
          for (forvar310 = (1'h0); (forvar310 < (2'h2)); forvar310 = (forvar310 + (1'h1)))
            begin
              reg311 <= (+(~&$signed(((~reg307) ?
                  (reg299 ? reg302 : wire295) : {wire298, reg299}))));
              reg312 <= ({(~^(^~$signed(forvar310)))} ?
                  $unsigned(reg305) : reg306);
              reg313 <= reg311;
              reg314 <= (&wire297);
              reg315 <= reg302[(2'h3):(2'h2)];
            end
        end
      for (forvar316 = (1'h0); (forvar316 < (3'h4)); forvar316 = (forvar316 + (1'h1)))
        begin
          reg317 <= reg301[(3'h6):(1'h0)];
          reg318 = ((($unsigned({reg301}) ?
              reg308 : wire298) == (wire296[(5'h12):(5'h11)] ^~ (^$signed(reg306)))) <= reg304[(4'h9):(1'h0)]);
        end
      reg319 <= wire297[(3'h6):(3'h6)];
    end
  always
    @(posedge clk) begin
      reg320 = $unsigned((&(|$unsigned((wire295 ? reg303 : reg319)))));
    end
  always
    @(posedge clk) begin
      for (forvar321 = (1'h0); (forvar321 < (2'h3)); forvar321 = (forvar321 + (1'h1)))
        begin
          reg322 <= (($signed({$signed(reg312), (~|reg301)}) ?
              (($signed(reg315) == (wire298 * reg308)) ?
                  ({reg317, reg300} ?
                      $unsigned(reg299) : wire297) : ((8'hac) == (wire296 ?
                      reg313 : reg315))) : $unsigned((|$unsigned(reg305)))) >= (reg305[(4'ha):(3'h5)] ^ $unsigned((wire298[(1'h1):(1'h0)] ?
              (^reg313) : (reg303 >> reg314)))));
        end
      reg323 <= (reg319[(5'h13):(4'hd)] ?
          $signed(($unsigned(reg319[(3'h4):(3'h4)]) ?
              $signed($signed((8'hbb))) : ($unsigned(reg312) ?
                  $unsigned(wire298) : wire296))) : ($signed(reg304) <= {$unsigned(reg313[(1'h0):(1'h0)])}));
      reg324 <= (|((reg305[(2'h3):(1'h1)] <<< wire297[(2'h2):(1'h1)]) ?
          $unsigned($signed(reg322[(3'h4):(1'h1)])) : ({$signed((8'hb7)),
                  (reg319 ^ reg307)} ?
              (reg299[(4'hb):(4'h8)] ^ (8'ha3)) : reg314[(1'h0):(1'h0)])));
    end
  assign wire325 = $unsigned(wire297);
  always
    @(posedge clk) begin
      for (forvar326 = (1'h0); (forvar326 < (1'h0)); forvar326 = (forvar326 + (1'h1)))
        begin
          reg327 <= $signed((~&$unsigned($unsigned($signed(reg301)))));
        end
      reg328 <= {(8'hbe)};
      if ($unsigned(forvar326[(3'h7):(2'h3)]))
        begin
          reg329 = (-$unsigned({$signed(forvar326)}));
          reg330 <= (((^~reg313) ~^ reg322[(2'h2):(1'h1)]) >> $unsigned(reg315[(1'h1):(1'h1)]));
        end
      else
        begin
          reg329 = reg306[(4'h9):(2'h2)];
        end
      reg331 <= $signed(wire298[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg332 <= wire295[(3'h6):(1'h0)];
      reg333 = $unsigned(wire296[(1'h0):(1'h0)]);
      reg334 <= {$signed($unsigned(((reg308 ? reg308 : reg313) ?
              (~|(8'ha6)) : reg315[(1'h0):(1'h0)]))),
          $unsigned(reg313)};
      reg335 <= (~|reg330);
    end
  assign wire336 = reg323;
  assign wire337 = (~{$unsigned(reg335[(3'h5):(1'h1)])});
  assign wire338 = $unsigned((&(($unsigned((8'hbb)) ?
                       (wire297 ?
                           reg328 : wire337) : reg335[(2'h2):(2'h2)]) <= $signed(wire336[(1'h1):(1'h1)]))));
  always
    @(posedge clk) begin
      reg339 <= (!$signed($unsigned($signed($unsigned(reg324)))));
      reg340 <= reg332;
      reg341 <= (-reg327[(3'h5):(3'h4)]);
      if (((reg327[(2'h3):(1'h0)] ?
              (-reg322) : $signed($signed($signed(reg301)))) ?
          {$signed((8'hb6))} : reg335[(3'h4):(2'h2)]))
        begin
          reg342 <= $signed((&{$signed($unsigned(reg307)),
              (~|$unsigned(reg311))}));
          reg343 <= (-$unsigned($signed(wire298[(1'h0):(1'h0)])));
        end
      else
        begin
          reg342 <= $signed((wire297 ?
              (reg299 ?
                  reg317[(2'h3):(2'h2)] : ((reg313 ? reg331 : reg340) ?
                      $signed(wire336) : $signed(reg313))) : reg315));
        end
      if (((reg308 >>> ((reg308[(2'h2):(1'h1)] != reg303) >>> reg304[(1'h0):(1'h0)])) ?
          $unsigned(wire298[(1'h1):(1'h1)]) : (-$unsigned(reg312[(3'h6):(2'h2)]))))
        begin
          for (forvar344 = (1'h0); (forvar344 < (1'h0)); forvar344 = (forvar344 + (1'h1)))
            begin
              reg345 <= ((~|((&reg315[(1'h1):(1'h0)]) ?
                  (8'ha9) : (reg342 == ((8'hb4) ?
                      reg313 : reg306)))) ~^ (((~|(reg311 ^~ reg301)) ?
                  (~reg301[(1'h0):(1'h0)]) : (8'ha7)) == (~&(^reg300[(1'h0):(1'h0)]))));
              reg346 <= ((($signed((|reg328)) > $signed((reg302 ?
                  reg319 : wire336))) | ($signed(reg335[(1'h1):(1'h1)]) <= $signed((~^reg324)))) ^~ (~&wire298));
              reg347 <= ($signed($signed({(!(8'h9e)),
                  $signed((8'hbf))})) * ((reg339 ?
                      ($unsigned((8'ha6)) ?
                          reg303 : reg324[(3'h5):(3'h4)]) : (reg342 ?
                          (reg346 ?
                              (7'h41) : reg323) : reg313[(5'h15):(4'hc)])) ?
                  $signed((reg341 ~^ $signed(reg340))) : $signed(wire298)));
              reg348 <= $signed(((&$unsigned((8'h9e))) != reg314));
            end
          reg349 <= (8'ha2);
        end
      else
        begin
          reg344 <= (~|(&wire296[(4'hc):(3'h7)]));
          reg345 <= (wire298[(1'h0):(1'h0)] ?
              {reg311} : (&(+{(8'hba), $unsigned(reg346)})));
        end
    end
  always
    @(posedge clk) begin
      reg350 <= wire325;
      reg351 <= $signed($unsigned($unsigned($unsigned($signed(wire297)))));
    end
  always
    @(posedge clk) begin
      for (forvar352 = (1'h0); (forvar352 < (2'h3)); forvar352 = (forvar352 + (1'h1)))
        begin
          reg353 <= ((~reg350[(2'h3):(1'h1)]) > (+$signed($unsigned((~&reg308)))));
          reg354 <= (^reg323);
          reg355 <= reg340[(4'h9):(3'h5)];
          reg356 <= reg339[(4'h9):(4'h9)];
          reg357 <= $signed($unsigned(wire298[(1'h1):(1'h0)]));
        end
      reg358 <= $unsigned($signed(reg347[(3'h4):(1'h0)]));
      reg359 <= reg331[(5'h11):(5'h10)];
    end
  assign wire360 = wire296;
  always
    @(posedge clk) begin
      for (forvar361 = (1'h0); (forvar361 < (1'h0)); forvar361 = (forvar361 + (1'h1)))
        begin
          reg362 <= (reg319[(2'h2):(1'h1)] && reg311);
          if (reg305)
            begin
              reg363 <= (^($unsigned((!(!reg348))) ?
                  $unsigned(((reg307 <<< reg359) | reg313)) : $unsigned((|(&reg302)))));
            end
          else
            begin
              reg363 <= $signed((8'ha2));
              reg364 = reg313[(3'h5):(1'h0)];
              reg365 <= wire336;
              reg366 = $signed(reg315[(1'h0):(1'h0)]);
              reg367 <= $signed(((|$signed($signed(reg303))) ~^ ({$unsigned(reg304)} >>> ((~|wire360) ?
                  (reg305 == (8'ha1)) : $unsigned(reg331)))));
            end
          if ((reg302 >= (!(reg315[(1'h0):(1'h0)] ?
              $signed((~^reg314)) : (((8'ha0) ? wire296 : (8'ha7)) ?
                  $signed(reg344) : (+forvar361))))))
            begin
              reg368 <= $unsigned((((~|(~&reg317)) < $unsigned((reg362 >> reg327))) ?
                  ($signed($signed(reg339)) ?
                      reg300 : reg306) : $unsigned({forvar361[(1'h1):(1'h0)]})));
              reg369 <= (~|((^~($unsigned((8'hbb)) && wire338)) <= forvar361[(4'hd):(4'h9)]));
              reg370 = (-(+{((reg301 ^ forvar361) <<< reg301),
                  $unsigned($signed((8'h9c)))}));
              reg371 <= ((7'h44) ? wire325 : (&$signed(reg343)));
              reg372 <= $unsigned(reg299);
            end
          else
            begin
              reg368 <= reg356;
              reg369 <= ({((|(reg302 ? reg307 : (8'hbd))) ?
                      ($signed(reg343) >= (reg301 ?
                          wire296 : reg349)) : reg304[(4'h9):(4'h8)]),
                  reg330} <<< (($signed({reg324}) ?
                      reg349 : (reg364[(4'hf):(3'h5)] > reg349)) ?
                  wire296 : reg367));
              reg371 <= (~&reg365);
            end
          reg373 <= (^reg306[(1'h0):(1'h0)]);
        end
    end
  always
    @(posedge clk) begin
      reg374 <= $unsigned(reg330);
      reg375 <= (((((reg317 - reg358) << (reg311 ? (8'hbc) : reg371)) ?
          (^~$unsigned(reg359)) : $unsigned(wire298[(1'h1):(1'h1)])) ~^ $signed($unsigned((^~reg323)))) + $signed($unsigned(($unsigned(reg355) ^~ reg308))));
      reg376 <= $signed((reg343 ?
          wire295[(2'h3):(2'h2)] : (~^($unsigned((8'haf)) + $signed(reg340)))));
      if (((($unsigned((reg350 ? reg362 : reg363)) ?
                  reg368[(2'h2):(1'h1)] : ((reg359 ? wire325 : reg327) ?
                      (reg357 ? reg300 : reg351) : (|reg351))) ?
              reg335[(1'h1):(1'h1)] : (8'h9c)) ?
          (~$unsigned({((8'hba) ?
                  (8'haa) : (8'ha0))})) : (wire295 | ($signed($unsigned(reg303)) ?
              {reg323[(5'h11):(2'h3)], (&(8'ha8))} : $unsigned((reg330 ?
                  (8'ha0) : wire360))))))
        begin
          reg377 <= reg369;
          reg378 <= reg332[(2'h2):(2'h2)];
          reg379 <= (reg319 ?
              (+reg367[(3'h5):(2'h3)]) : ($signed(($unsigned(reg371) || (~&wire297))) > $signed(reg304)));
          for (forvar380 = (1'h0); (forvar380 < (3'h4)); forvar380 = (forvar380 + (1'h1)))
            begin
              reg381 <= (((~{(reg319 | (8'hb5))}) ?
                  (reg362[(2'h2):(2'h2)] ?
                      reg305 : $unsigned(wire338)) : ($unsigned((reg308 >> reg356)) | ((~wire297) & $unsigned(reg307)))) + $signed({{$signed(wire337)}}));
              reg382 <= reg302[(2'h2):(1'h1)];
              reg383 <= ({({reg376[(4'ha):(4'h8)], (^~reg307)} ?
                      reg312[(3'h6):(2'h2)] : $unsigned(reg335[(2'h2):(2'h2)]))} | $unsigned(wire360));
            end
          reg384 <= $signed((((((8'hb3) & reg304) ?
                  (forvar380 >> reg369) : (reg373 ? reg363 : reg362)) ?
              (forvar380 >>> reg302[(4'h8):(4'h8)]) : (reg315 >= (reg368 ?
                  (8'haf) : reg300))) & reg372[(1'h1):(1'h1)]));
        end
      else
        begin
          reg377 <= $signed((!$signed($unsigned((&reg314)))));
        end
    end
  assign wire385 = ((~&((&reg340[(5'h12):(2'h2)]) ^ ({reg342, reg351} ?
                       ((8'hb7) >= reg379) : (reg300 ?
                           wire337 : wire295)))) - $signed((~^$signed($signed(reg365)))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module145  (y, clk, wire149, wire148, wire147, wire146);
  output wire [(32'h746):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hb):(1'h0)] wire149;
  input wire [(5'h14):(1'h0)] wire148;
  input wire [(4'hd):(1'h0)] wire147;
  input wire signed [(5'h12):(1'h0)] wire146;
  wire [(4'h8):(1'h0)] wire256;
  wire signed [(4'h9):(1'h0)] wire197;
  wire signed [(3'h4):(1'h0)] wire196;
  wire [(5'h15):(1'h0)] wire195;
  wire signed [(3'h6):(1'h0)] wire194;
  wire [(5'h10):(1'h0)] wire193;
  wire [(3'h7):(1'h0)] wire179;
  wire [(3'h4):(1'h0)] wire178;
  wire [(4'hb):(1'h0)] wire156;
  wire [(5'h12):(1'h0)] wire151;
  wire [(4'he):(1'h0)] wire150;
  reg [(4'he):(1'h0)] reg288 = (1'h0);
  reg [(4'h8):(1'h0)] reg286 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg284 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg283 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg281 = (1'h0);
  reg [(4'h8):(1'h0)] reg280 = (1'h0);
  reg [(5'h11):(1'h0)] reg279 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg278 = (1'h0);
  reg [(5'h14):(1'h0)] reg276 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg274 = (1'h0);
  reg [(5'h12):(1'h0)] reg272 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg270 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg269 = (1'h0);
  reg [(5'h11):(1'h0)] reg265 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg261 = (1'h0);
  reg [(4'h8):(1'h0)] reg260 = (1'h0);
  reg [(4'hc):(1'h0)] reg258 = (1'h0);
  reg [(5'h15):(1'h0)] reg257 = (1'h0);
  reg [(4'hd):(1'h0)] reg255 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg254 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg253 = (1'h0);
  reg [(4'hd):(1'h0)] reg252 = (1'h0);
  reg [(5'h14):(1'h0)] reg251 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg250 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg249 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg247 = (1'h0);
  reg [(4'he):(1'h0)] reg246 = (1'h0);
  reg [(4'hd):(1'h0)] reg245 = (1'h0);
  reg [(5'h11):(1'h0)] reg244 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg243 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg242 = (1'h0);
  reg [(3'h6):(1'h0)] reg241 = (1'h0);
  reg [(4'hf):(1'h0)] reg239 = (1'h0);
  reg [(4'hf):(1'h0)] reg238 = (1'h0);
  reg [(5'h13):(1'h0)] reg237 = (1'h0);
  reg [(4'hd):(1'h0)] reg230 = (1'h0);
  reg signed [(4'he):(1'h0)] reg235 = (1'h0);
  reg [(3'h7):(1'h0)] reg234 = (1'h0);
  reg [(5'h12):(1'h0)] reg233 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg231 = (1'h0);
  reg [(4'ha):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg228 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg225 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg224 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg223 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg221 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg217 = (1'h0);
  reg [(4'h9):(1'h0)] reg216 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg198 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg215 = (1'h0);
  reg [(4'he):(1'h0)] reg214 = (1'h0);
  reg [(5'h12):(1'h0)] reg213 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg212 = (1'h0);
  reg signed [(4'he):(1'h0)] reg211 = (1'h0);
  reg [(4'he):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg208 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg207 = (1'h0);
  reg [(4'hf):(1'h0)] reg206 = (1'h0);
  reg [(4'ha):(1'h0)] reg205 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg203 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg201 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg200 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg199 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg192 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg191 = (1'h0);
  reg [(5'h12):(1'h0)] reg184 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg190 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg189 = (1'h0);
  reg [(4'hc):(1'h0)] reg188 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg187 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg186 = (1'h0);
  reg [(4'hd):(1'h0)] reg182 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg177 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg176 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg175 = (1'h0);
  reg [(4'hc):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg173 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg171 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg170 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg168 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg167 = (1'h0);
  reg [(5'h11):(1'h0)] reg166 = (1'h0);
  reg [(4'h8):(1'h0)] reg165 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg162 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg161 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg160 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg157 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg155 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg154 = (1'h0);
  reg [(3'h4):(1'h0)] reg153 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg152 = (1'h0);
  reg [(5'h13):(1'h0)] reg289 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg287 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg285 = (1'h0);
  reg [(4'ha):(1'h0)] reg282 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg277 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar275 = (1'h0);
  reg [(5'h13):(1'h0)] forvar273 = (1'h0);
  reg [(4'hf):(1'h0)] forvar271 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg268 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg267 = (1'h0);
  reg [(4'h9):(1'h0)] forvar266 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg264 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg262 = (1'h0);
  reg [(5'h12):(1'h0)] reg259 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg248 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar240 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg236 = (1'h0);
  reg [(5'h14):(1'h0)] forvar230 = (1'h0);
  reg signed [(4'he):(1'h0)] reg227 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg219 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar210 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar198 = (1'h0);
  reg [(4'he):(1'h0)] reg185 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar184 = (1'h0);
  reg [(5'h11):(1'h0)] reg183 = (1'h0);
  reg [(4'ha):(1'h0)] reg181 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg180 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg169 = (1'h0);
  reg [(4'he):(1'h0)] reg172 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar169 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg164 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar163 = (1'h0);
  reg [(5'h10):(1'h0)] forvar158 = (1'h0);
  assign y = {wire256,
                 wire197,
                 wire196,
                 wire195,
                 wire194,
                 wire193,
                 wire179,
                 wire178,
                 wire156,
                 wire151,
                 wire150,
                 reg288,
                 reg286,
                 reg284,
                 reg283,
                 reg281,
                 reg280,
                 reg279,
                 reg278,
                 reg276,
                 reg274,
                 reg272,
                 reg270,
                 reg269,
                 reg265,
                 reg263,
                 reg261,
                 reg260,
                 reg258,
                 reg257,
                 reg255,
                 reg254,
                 reg253,
                 reg252,
                 reg251,
                 reg250,
                 reg249,
                 reg247,
                 reg246,
                 reg245,
                 reg244,
                 reg243,
                 reg242,
                 reg241,
                 reg239,
                 reg238,
                 reg237,
                 reg230,
                 reg235,
                 reg234,
                 reg233,
                 reg232,
                 reg231,
                 reg229,
                 reg228,
                 reg226,
                 reg225,
                 reg224,
                 reg223,
                 reg222,
                 reg221,
                 reg220,
                 reg218,
                 reg217,
                 reg216,
                 reg198,
                 reg215,
                 reg214,
                 reg213,
                 reg212,
                 reg211,
                 reg209,
                 reg208,
                 reg207,
                 reg206,
                 reg205,
                 reg204,
                 reg203,
                 reg202,
                 reg201,
                 reg200,
                 reg199,
                 reg192,
                 reg191,
                 reg184,
                 reg190,
                 reg189,
                 reg188,
                 reg187,
                 reg186,
                 reg182,
                 reg177,
                 reg176,
                 reg175,
                 reg174,
                 reg173,
                 reg171,
                 reg170,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg162,
                 reg161,
                 reg160,
                 reg159,
                 reg157,
                 reg155,
                 reg154,
                 reg153,
                 reg152,
                 reg289,
                 reg287,
                 reg285,
                 reg282,
                 reg277,
                 forvar275,
                 forvar273,
                 forvar271,
                 reg268,
                 reg267,
                 forvar266,
                 reg264,
                 reg262,
                 reg259,
                 reg248,
                 forvar240,
                 reg236,
                 forvar230,
                 reg227,
                 reg219,
                 forvar210,
                 forvar198,
                 reg185,
                 forvar184,
                 reg183,
                 reg181,
                 reg180,
                 reg169,
                 reg172,
                 forvar169,
                 reg164,
                 forvar163,
                 forvar158,
                 (1'h0)};
  assign wire150 = $signed((wire147[(1'h1):(1'h1)] ?
                       (wire148[(5'h10):(1'h1)] ~^ (wire147 <<< wire147[(3'h6):(3'h4)])) : wire149));
  assign wire151 = ({$signed($signed((wire146 ^~ wire149))), wire147} ?
                       ($unsigned((&wire147)) | wire150[(4'hb):(4'hb)]) : wire148);
  always
    @(posedge clk) begin
      reg152 <= (+wire151[(2'h2):(1'h1)]);
      reg153 <= {(!(&wire150)),
          (($unsigned($unsigned(wire146)) ?
              ($signed(reg152) ?
                  (+wire148) : (~wire148)) : reg152) != wire151[(5'h10):(5'h10)])};
      reg154 <= wire146;
      reg155 <= (wire150[(4'hd):(4'hc)] ? wire147 : $unsigned(wire150));
    end
  assign wire156 = $signed(({$unsigned(wire146)} ?
                       wire146[(2'h3):(1'h1)] : (reg155 ?
                           $unsigned(reg153) : wire150)));
  always
    @(posedge clk) begin
      reg157 <= $signed((~|(^reg152)));
      for (forvar158 = (1'h0); (forvar158 < (3'h4)); forvar158 = (forvar158 + (1'h1)))
        begin
          reg159 <= reg152;
          reg160 <= {($unsigned($signed((^~wire147))) >>> wire148),
              $unsigned((forvar158[(4'hf):(4'hb)] * (~^((8'haf) ?
                  wire150 : reg155))))};
          if ($unsigned($unsigned(((~|$signed(wire151)) ?
              {wire151} : (~reg154)))))
            begin
              reg161 <= reg153[(2'h2):(2'h2)];
              reg162 <= ($signed(((~wire156) ?
                      wire150[(4'ha):(4'ha)] : reg161)) ?
                  (wire150[(1'h0):(1'h0)] ?
                      (^~(-wire151[(3'h4):(1'h0)])) : wire151[(3'h6):(3'h6)]) : $unsigned($signed(reg153[(2'h2):(2'h2)])));
            end
          else
            begin
              reg161 <= reg152[(4'ha):(4'h8)];
              reg162 <= {reg157,
                  $signed(($unsigned(wire156[(3'h4):(1'h1)]) ?
                      (-(reg153 ?
                          wire147 : wire149)) : wire149[(2'h3):(2'h2)]))};
            end
          for (forvar163 = (1'h0); (forvar163 < (2'h2)); forvar163 = (forvar163 + (1'h1)))
            begin
              reg164 = {reg161, (7'h40)};
              reg165 <= reg164;
            end
        end
      reg166 <= (8'ha6);
      if ($unsigned((($unsigned($unsigned((8'hba))) <<< ((^~(8'ha5)) ?
          {wire156} : reg154[(3'h6):(2'h2)])) & wire156)))
        begin
          reg167 <= $unsigned({(^~wire156[(3'h6):(3'h4)]),
              wire150[(4'hd):(1'h1)]});
          reg168 <= wire149;
          for (forvar169 = (1'h0); (forvar169 < (1'h0)); forvar169 = (forvar169 + (1'h1)))
            begin
              reg170 <= (reg164 >>> (~|(~(reg166[(2'h3):(1'h0)] ?
                  (reg162 ~^ forvar163) : (reg161 & reg155)))));
              reg171 <= {wire151[(3'h5):(3'h4)]};
              reg172 = ($unsigned(wire147) != wire147[(3'h5):(3'h5)]);
            end
        end
      else
        begin
          if ((^$signed(((reg155[(2'h2):(1'h1)] <= (reg168 ?
              wire149 : forvar163)) ~^ (+$signed(wire156))))))
            begin
              reg167 <= reg162[(1'h1):(1'h0)];
              reg168 <= (~$unsigned(($signed(reg164[(1'h0):(1'h0)]) - ($signed(reg155) ?
                  (|(8'hae)) : $unsigned(reg152)))));
              reg169 = $signed((8'ha0));
              reg170 <= (8'hac);
            end
          else
            begin
              reg167 <= {{reg159[(3'h4):(1'h1)], reg152[(4'ha):(1'h0)]}};
              reg168 <= ($signed(($unsigned(wire150[(1'h0):(1'h0)]) >= reg165[(4'h8):(1'h1)])) ?
                  $signed(((^~(8'hb6)) ?
                      {$unsigned((8'hb4)),
                          reg168[(3'h7):(3'h5)]} : reg170[(2'h2):(2'h2)])) : $unsigned((-wire149)));
            end
        end
      reg173 <= $unsigned(reg165[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg174 <= (~(^~($unsigned({reg166}) ?
          $signed((wire147 + wire156)) : {$unsigned((8'hb3)),
              ((8'hbf) ~^ wire148)})));
      reg175 <= ((8'hb0) * $unsigned(((wire149[(2'h3):(2'h3)] ?
              $unsigned(reg173) : $unsigned(reg167)) ?
          $unsigned(reg152[(4'h8):(4'h8)]) : (|(&reg159)))));
      reg176 <= wire148[(3'h5):(2'h3)];
      reg177 <= $signed($signed(reg176[(3'h5):(3'h4)]));
    end
  assign wire178 = (|{($signed(wire156) >> {(wire150 && reg166),
                           $unsigned(wire147)})});
  assign wire179 = reg176[(5'h13):(2'h3)];
  always
    @(posedge clk) begin
      reg180 = wire178;
      if ($signed(((({reg171} * $signed(reg171)) ?
              ((8'hab) == $signed(reg165)) : (+reg170)) ?
          {(reg157[(5'h13):(2'h2)] ?
                  reg177[(4'h8):(2'h2)] : $unsigned((8'hb2))),
              ($unsigned(reg170) ?
                  (wire178 ~^ reg152) : $unsigned(reg168))} : (&$signed((reg161 ?
              reg161 : reg155))))))
        begin
          reg181 = (((&wire151) >>> (~{reg165[(3'h4):(3'h4)],
              (^reg167)})) & $unsigned(reg162));
          reg182 <= (reg170 <= $signed(reg177));
          reg183 = ($unsigned(reg152[(3'h5):(2'h3)]) ?
              $unsigned($signed($signed((|reg153)))) : wire148[(1'h1):(1'h1)]);
          for (forvar184 = (1'h0); (forvar184 < (2'h3)); forvar184 = (forvar184 + (1'h1)))
            begin
              reg185 = (+wire147);
              reg186 <= $signed($unsigned(reg160));
              reg187 <= {$signed(($unsigned({reg152, (8'hb7)}) ?
                      (((8'ha8) >>> reg171) ?
                          wire156 : (reg186 ?
                              reg186 : (8'h9e))) : $signed((~&reg186)))),
                  wire178[(1'h0):(1'h0)]};
              reg188 <= (^~(~$unsigned((~^$unsigned(forvar184)))));
              reg189 <= $unsigned(wire147[(4'hc):(4'h8)]);
            end
          reg190 <= reg183;
        end
      else
        begin
          reg182 <= wire148[(4'h8):(3'h5)];
          reg184 <= (reg161 ?
              ((($unsigned(reg171) ? (~reg154) : (reg185 <= wire179)) ?
                  $signed(forvar184) : (wire148[(5'h12):(4'he)] ?
                      reg153[(1'h1):(1'h1)] : (reg154 ?
                          (8'had) : reg180))) << $unsigned({$signed(reg171)})) : ($unsigned((((8'hbd) ?
                      reg161 : reg153) ?
                  (reg171 > reg160) : reg189)) == reg166));
          reg186 <= ((reg175 ? (^reg187) : reg182) >= reg157);
          if ((!$unsigned({wire147[(4'ha):(3'h5)]})))
            begin
              reg187 <= $signed({reg184[(4'hb):(4'ha)]});
            end
          else
            begin
              reg187 <= (~|({$unsigned((reg188 ? reg190 : (8'h9e))),
                      (^(reg181 || reg165))} ?
                  reg174 : wire179));
            end
          if ($unsigned(reg153[(3'h4):(2'h3)]))
            begin
              reg188 <= (^~$signed(($signed(wire156[(1'h0):(1'h0)]) ?
                  (7'h40) : wire146)));
              reg189 <= (({((forvar184 >> reg184) ?
                          reg171 : wire150[(4'he):(3'h5)])} <= $unsigned(wire156[(3'h5):(3'h4)])) ?
                  reg174[(3'h4):(2'h2)] : (~&$unsigned(reg171[(3'h5):(3'h5)])));
            end
          else
            begin
              reg188 <= {reg174};
              reg189 <= (((~|$unsigned(reg181[(2'h2):(2'h2)])) << ({(reg166 >>> reg190)} ?
                      reg174[(4'h8):(1'h1)] : (+{reg168, reg186}))) ?
                  (^reg186[(3'h7):(2'h3)]) : $signed($unsigned(reg161[(3'h7):(3'h6)])));
            end
        end
      reg191 <= $unsigned($signed((^reg165[(1'h0):(1'h0)])));
      reg192 <= {($unsigned(reg171[(4'h8):(1'h0)]) ~^ ($unsigned(reg167[(1'h1):(1'h0)]) <<< {reg153[(2'h2):(1'h1)]})),
          wire146};
    end
  assign wire193 = (reg192 ?
                       (8'hbf) : $signed(($unsigned($unsigned(reg159)) || reg168)));
  assign wire194 = ((|$signed($signed((^~reg192)))) ?
                       (reg182 >> ((-(^~(8'hb6))) ?
                           {(reg174 ? reg157 : (8'haf)),
                               wire193[(4'ha):(4'h8)]} : {(wire178 < reg191)})) : $signed(reg161));
  assign wire195 = ({reg170} != $unsigned((~&$unsigned($unsigned(reg177)))));
  assign wire196 = $signed((((8'ha8) ?
                       $signed((reg174 ?
                           reg152 : reg157)) : wire178) * (+reg162[(2'h3):(1'h1)])));
  assign wire197 = wire194[(3'h6):(3'h6)];
  always
    @(posedge clk) begin
      if (((($unsigned({reg157}) ? (8'hb3) : $unsigned((&reg171))) ?
              reg184 : ((~&$unsigned((8'hb8))) ?
                  $unsigned((reg152 ?
                      wire178 : reg168)) : $unsigned($unsigned(reg187)))) ?
          ((~^($unsigned(reg166) || (reg165 ? reg186 : reg186))) ?
              $signed((wire179 ^~ (wire178 - (7'h43)))) : (($unsigned(reg162) ^ reg174) ?
                  ($signed((8'hbc)) ?
                      (reg177 + reg152) : {(8'hb0), (8'ha1)}) : {(wire194 ?
                          (8'h9d) : wire156),
                      $signed(reg182)})) : reg161))
        begin
          for (forvar198 = (1'h0); (forvar198 < (1'h0)); forvar198 = (forvar198 + (1'h1)))
            begin
              reg199 <= (($signed((reg175 ?
                      (!wire178) : reg182[(4'h9):(3'h7)])) < (!$signed(reg159[(1'h0):(1'h0)]))) ?
                  (^~(^$unsigned(((8'hae) + reg159)))) : {$unsigned(reg167[(3'h4):(1'h1)]),
                      reg189});
              reg200 <= reg192[(2'h2):(2'h2)];
              reg201 <= (wire178 >> forvar198[(2'h2):(1'h0)]);
              reg202 <= (reg184[(5'h11):(3'h4)] ?
                  (|{(reg173 ?
                          (reg159 >> wire193) : $unsigned(reg188))}) : (8'hb5));
              reg203 <= (($unsigned($unsigned($signed(wire150))) ^~ reg159[(3'h5):(2'h2)]) >= (8'haa));
            end
          reg204 <= reg186;
          if ($signed(($unsigned((((8'ha7) ?
                  reg173 : wire149) < wire179[(3'h7):(3'h6)])) ?
              $signed($signed({wire151})) : (!(&$signed(reg199))))))
            begin
              reg205 <= (^(~^reg191[(1'h0):(1'h0)]));
              reg206 <= (reg154 >>> (reg186[(3'h4):(1'h0)] ~^ ($signed((~&reg200)) >= reg159[(3'h5):(1'h0)])));
              reg207 <= (((~^(^reg187)) ?
                  (($unsigned((8'hb0)) >= (reg205 <<< wire193)) + reg155) : (reg176[(1'h1):(1'h1)] ?
                      wire148[(4'hb):(3'h7)] : $unsigned((reg176 >> wire149)))) < {($unsigned($signed(reg184)) ?
                      ((~|reg204) ?
                          reg177[(4'ha):(3'h5)] : $signed(reg204)) : ((reg173 | reg167) ?
                          (reg155 != reg203) : $unsigned(reg177))),
                  (+($unsigned(reg188) ?
                      reg153[(1'h0):(1'h0)] : (reg165 >= forvar198)))});
              reg208 <= {{(~^reg186[(1'h0):(1'h0)]),
                      $unsigned((((8'h9e) << reg154) ?
                          reg184 : $signed(wire149)))}};
            end
          else
            begin
              reg205 <= (((wire148[(1'h1):(1'h0)] & (reg175[(4'hb):(1'h0)] ?
                      {(8'hb9)} : (reg167 ? reg168 : wire179))) ?
                  {reg155[(3'h5):(1'h0)]} : $unsigned(((wire156 | wire197) ?
                      {reg203, reg174} : (reg202 ?
                          wire148 : (8'ha7))))) & $unsigned(reg175[(3'h7):(3'h6)]));
            end
          reg209 <= ($signed((($signed(reg182) == $signed(reg173)) && (+reg177))) ?
              {(~&($unsigned((8'ha0)) != (reg153 ?
                      reg174 : reg189)))} : {(&((~^reg187) ?
                      (wire178 ? reg184 : reg205) : $signed(reg204))),
                  ({(~&reg168), $unsigned(reg167)} ?
                      ((!reg174) <<< $signed((8'hb1))) : $unsigned(reg166[(2'h3):(2'h2)]))});
          for (forvar210 = (1'h0); (forvar210 < (2'h3)); forvar210 = (forvar210 + (1'h1)))
            begin
              reg211 <= reg189;
              reg212 <= $signed((!(&{(reg186 ? wire147 : wire196),
                  $unsigned(reg209)})));
              reg213 <= {$signed(($unsigned((reg152 - reg161)) ?
                      reg187 : reg211[(4'h9):(1'h1)])),
                  (+reg199)};
              reg214 <= wire194[(3'h4):(1'h1)];
              reg215 <= $unsigned((((reg203[(3'h6):(1'h1)] ^ (wire150 ?
                      wire178 : wire151)) >> $signed((reg189 && reg189))) ?
                  {{{wire156, forvar198},
                          (reg207 * reg212)}} : $unsigned(((wire179 - reg168) && $unsigned(reg160)))));
            end
        end
      else
        begin
          reg198 <= $unsigned(reg174[(4'hc):(2'h2)]);
        end
      if ($unsigned($signed(((reg160 ? {reg213} : (reg199 == (8'hbc))) ?
          wire150 : $signed($unsigned(reg175))))))
        begin
          reg216 <= (&(~&(~reg192)));
          reg217 <= $signed((|(reg198[(1'h0):(1'h0)] > $signed(reg165))));
        end
      else
        begin
          reg216 <= (~|$signed(reg188));
        end
      reg218 <= (~|wire149[(4'hb):(2'h3)]);
      reg219 = ({$signed({{reg207, reg173}, (~|(8'ha1))}),
              {((+reg198) ? $signed(wire147) : $unsigned(reg176))}} ?
          reg184 : (wire151[(1'h1):(1'h0)] <= ((|(reg159 ?
              reg173 : reg215)) ^ {(-reg162), $signed(reg218)})));
    end
  always
    @(posedge clk) begin
      reg220 <= ({$signed(reg200[(2'h2):(1'h1)])} ^~ $signed(reg201[(4'h9):(1'h0)]));
      reg221 <= reg159[(4'h8):(1'h1)];
      reg222 <= {$signed($signed({(reg211 ? wire195 : reg217)}))};
      reg223 <= reg189;
      reg224 <= $unsigned((-reg187[(2'h2):(2'h2)]));
    end
  always
    @(posedge clk) begin
      if (($signed((8'hb7)) ?
          ($unsigned(((reg218 ?
              reg166 : reg203) >> (~&reg176))) ^ reg214) : reg174[(4'hc):(3'h6)]))
        begin
          if ((reg159[(4'h8):(1'h0)] & ({reg221,
              (~&(reg184 ?
                  reg177 : reg187))} & (~^$signed(reg218[(3'h5):(3'h4)])))))
            begin
              reg225 <= $signed(reg168[(3'h6):(1'h0)]);
              reg226 <= reg176;
              reg227 = $unsigned($signed({reg208, reg174}));
            end
          else
            begin
              reg225 <= $signed($unsigned((|reg174[(4'hb):(1'h0)])));
              reg226 <= reg215;
              reg228 <= (reg223[(4'hd):(4'hc)] || reg160[(1'h0):(1'h0)]);
              reg229 <= ($signed(reg176[(4'ha):(3'h6)]) ?
                  wire149 : reg174[(4'h8):(1'h1)]);
            end
          for (forvar230 = (1'h0); (forvar230 < (2'h3)); forvar230 = (forvar230 + (1'h1)))
            begin
              reg231 <= ($unsigned(reg160[(3'h6):(2'h3)]) && reg161);
              reg232 <= $signed((reg154[(1'h1):(1'h1)] ?
                  ((wire151 ? wire146[(4'he):(3'h5)] : (-(8'ha3))) ?
                      (^$unsigned(reg175)) : $signed($signed(reg207))) : wire149));
            end
          reg233 <= ((+reg161) * {(reg176[(3'h5):(2'h2)] != $signed(reg227))});
          reg234 <= (8'hbb);
          reg235 <= reg229[(1'h0):(1'h0)];
        end
      else
        begin
          reg225 <= reg228[(3'h7):(3'h4)];
          reg226 <= {$unsigned(reg157)};
          reg228 <= ($signed(reg206[(4'h9):(3'h5)]) >= (~($unsigned(reg209) ?
              $signed((~|reg189)) : ((reg204 ?
                  reg170 : wire147) ^~ (reg153 < wire151)))));
          if ((!({((^~(8'hbc)) ~^ (+reg155))} ^~ $signed(reg182[(4'h9):(4'h9)]))))
            begin
              reg229 <= (^~$unsigned((~^{reg213, $signed(wire146)})));
              reg230 <= $unsigned($signed({wire156}));
              reg231 <= reg168;
              reg232 <= (($unsigned($signed((reg162 + reg191))) ?
                  $unsigned(((reg199 ~^ reg231) ?
                      {reg232} : $unsigned((8'hae)))) : (reg155[(1'h1):(1'h0)] ?
                      (reg155[(3'h4):(1'h1)] + {reg228}) : (wire150[(3'h4):(1'h0)] ?
                          $unsigned((8'hb2)) : (reg234 ?
                              reg217 : reg173)))) ^~ ({((&reg182) ?
                          (reg173 || (8'haf)) : reg165[(2'h2):(2'h2)]),
                      ($signed(reg199) & (wire147 >= reg223))} ?
                  ($signed($signed((8'hae))) ?
                      $unsigned(reg235[(4'hc):(2'h3)]) : (+$unsigned(wire193))) : $unsigned(reg157)));
              reg233 <= reg175;
            end
          else
            begin
              reg229 <= $unsigned($unsigned(wire149[(1'h0):(1'h0)]));
              reg230 <= ($signed(reg168[(4'h8):(1'h0)]) & reg234);
              reg236 = reg154;
            end
          reg237 <= ($unsigned((reg206[(1'h0):(1'h0)] * (reg229[(3'h5):(3'h4)] && (reg201 << reg161)))) ?
              (^$signed(reg215)) : ($unsigned($unsigned($unsigned(reg236))) ?
                  (~&reg201[(5'h13):(3'h5)]) : $signed(((&forvar230) ?
                      (reg236 ? reg204 : reg232) : reg189[(4'ha):(4'ha)]))));
        end
      reg238 <= (reg223 || $signed($signed((((8'hb2) && wire156) ?
          (reg168 ? reg152 : reg209) : (reg223 ? reg188 : wire149)))));
      reg239 <= reg199;
    end
  always
    @(posedge clk) begin
      if ({$unsigned($unsigned((&{reg168}))),
          ($unsigned((~&reg199)) <= (~&($signed(reg166) ?
              ((8'ha0) ^ reg174) : $signed((8'haf)))))})
        begin
          for (forvar240 = (1'h0); (forvar240 < (3'h4)); forvar240 = (forvar240 + (1'h1)))
            begin
              reg241 <= $signed((reg220[(1'h0):(1'h0)] + $signed($signed($signed(reg176)))));
              reg242 <= reg187[(1'h0):(1'h0)];
              reg243 <= $signed(reg166);
              reg244 <= $unsigned(({$unsigned(reg199[(5'h10):(5'h10)])} << (~&reg223)));
              reg245 <= (-(reg182 >> reg182));
            end
          reg246 <= (~&$unsigned((((~|reg167) & reg209[(1'h0):(1'h0)]) ?
              {(~reg152), $unsigned(reg203)} : reg152[(2'h3):(2'h3)])));
          reg247 <= wire195;
        end
      else
        begin
          for (forvar240 = (1'h0); (forvar240 < (1'h0)); forvar240 = (forvar240 + (1'h1)))
            begin
              reg241 <= ((|(&reg160[(4'h8):(3'h7)])) < $unsigned(reg157));
              reg242 <= ((~^$signed($signed($unsigned(reg216)))) >> ((wire195[(4'hf):(3'h5)] ?
                  wire156[(3'h4):(3'h4)] : $unsigned(reg177)) ~^ reg175[(4'hd):(1'h0)]));
            end
          if ({($unsigned(((reg174 | reg239) <= (reg191 ? wire196 : reg159))) ?
                  (reg246[(1'h0):(1'h0)] | reg189) : $unsigned((reg162[(4'h8):(3'h4)] ?
                      reg243 : {reg205}))),
              wire149[(4'ha):(3'h4)]})
            begin
              reg243 <= {$signed((~$unsigned(reg222))), reg215};
              reg244 <= (reg199 ? reg205 : wire193);
            end
          else
            begin
              reg243 <= $unsigned((((|(~^reg190)) ^ {$signed(reg207)}) <<< reg224));
              reg244 <= ($unsigned(reg207) ?
                  reg201[(3'h5):(3'h5)] : $unsigned((wire146[(1'h0):(1'h0)] ?
                      {(+(8'ha7))} : ($unsigned(reg223) ?
                          (reg224 ? reg237 : reg229) : (^~(8'hae))))));
              reg245 <= reg235[(1'h1):(1'h1)];
            end
          reg248 = ((wire196 >> reg202[(2'h2):(1'h0)]) - (&reg191));
        end
      reg249 <= (reg200 ?
          reg168[(3'h6):(3'h6)] : ((reg217 ? reg168 : (8'hb0)) ?
              $unsigned((~&$signed(reg184))) : (&$unsigned((8'ha6)))));
      reg250 <= (+(reg238 ? reg173 : $unsigned(reg242)));
      reg251 <= $unsigned($signed($unsigned($signed(reg187))));
    end
  always
    @(posedge clk) begin
      reg252 <= (reg203 ?
          ((&$unsigned(((8'hb8) ?
              reg153 : wire193))) ~^ reg155[(1'h0):(1'h0)]) : (($unsigned($signed((8'ha6))) ?
              reg173 : reg215[(5'h10):(4'h9)]) >= reg221));
      reg253 <= $signed(reg177);
      reg254 <= (|(reg245[(2'h2):(1'h0)] * (reg243[(3'h6):(1'h1)] ?
          reg175 : (&(reg202 >> (8'hac))))));
      reg255 <= $signed(reg202);
    end
  assign wire256 = ($unsigned((8'hb4)) < (reg199 ^ $unsigned((reg215 == (reg247 >= reg242)))));
  always
    @(posedge clk) begin
      reg257 <= (~&reg177);
    end
  always
    @(posedge clk) begin
      if (reg154)
        begin
          reg258 <= (((^$unsigned((reg231 ? reg200 : (8'hb8)))) ?
              (reg247[(3'h4):(3'h4)] == reg244[(3'h7):(3'h6)]) : reg155[(1'h0):(1'h0)]) | {($signed((reg241 > wire149)) << (7'h42)),
              reg238});
        end
      else
        begin
          reg258 <= reg226[(1'h0):(1'h0)];
        end
      reg259 = $signed($signed((~&($unsigned((8'h9d)) <<< reg237[(4'hf):(4'hd)]))));
      if ((~|(~^$unsigned($unsigned(reg203)))))
        begin
          reg260 <= (~|({reg223} <= reg250[(2'h2):(2'h2)]));
          if (reg205)
            begin
              reg261 <= (~{$signed(reg171[(3'h5):(2'h2)])});
            end
          else
            begin
              reg262 = {reg216[(2'h3):(2'h2)], (^~reg202)};
              reg263 <= $signed(($signed({(reg220 < reg252),
                  wire178[(2'h2):(1'h0)]}) ^~ (((reg160 ?
                      reg222 : reg229) <<< (&reg230)) ?
                  {reg207} : reg253[(1'h0):(1'h0)])));
              reg264 = $signed(($signed((^(~^reg230))) < {{$signed(reg246),
                      $signed(reg250)},
                  reg251}));
            end
          reg265 <= {(-{((^(8'hb6)) - $unsigned(reg177))})};
          for (forvar266 = (1'h0); (forvar266 < (2'h2)); forvar266 = (forvar266 + (1'h1)))
            begin
              reg267 = {$unsigned(wire193)};
              reg268 = reg152;
            end
          reg269 <= $unsigned((~^$unsigned(((reg233 <= reg235) ?
              (reg202 << reg176) : wire195[(1'h0):(1'h0)]))));
        end
      else
        begin
          reg262 = reg214[(4'h9):(3'h5)];
          reg263 <= $signed((((reg255 ? (reg186 <= reg249) : wire156) ?
                  reg264 : (~|(reg184 ? reg241 : wire149))) ?
              reg202[(2'h3):(1'h0)] : $signed($signed((~|reg215)))));
        end
      reg270 <= $signed($unsigned(reg212));
      for (forvar271 = (1'h0); (forvar271 < (3'h4)); forvar271 = (forvar271 + (1'h1)))
        begin
          reg272 <= (!$signed($unsigned(({reg243} ?
              (reg220 ? (8'hb0) : reg214) : reg221[(4'h8):(1'h0)]))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar273 = (1'h0); (forvar273 < (3'h4)); forvar273 = (forvar273 + (1'h1)))
        begin
          reg274 <= reg162[(3'h4):(1'h0)];
          for (forvar275 = (1'h0); (forvar275 < (1'h0)); forvar275 = (forvar275 + (1'h1)))
            begin
              reg276 <= reg174;
              reg277 = (~wire193);
              reg278 <= (reg214[(3'h4):(2'h3)] ?
                  reg245[(1'h0):(1'h0)] : ((wire195[(4'he):(4'ha)] ?
                          (~^reg239) : reg263) ?
                      (reg214 + ($signed(reg253) < $signed(wire150))) : ($signed({(8'ha5)}) ?
                          ((reg229 & reg221) & reg176) : {(8'hbf)})));
              reg279 <= reg211[(4'hd):(4'h9)];
              reg280 <= (($signed((~&reg238[(3'h7):(3'h5)])) + $signed($unsigned(reg217[(4'he):(4'hc)]))) <<< (^$unsigned({(^~wire196)})));
            end
          reg281 <= ({(^{(+(7'h41))}),
              ((reg217 ?
                  (reg182 > reg280) : $unsigned(reg233)) < reg191[(1'h0):(1'h0)])} >= ((&(~^{reg265})) ?
              {wire193, reg187} : (^$unsigned(((8'hbf) + reg155)))));
          reg282 = ({((reg187[(2'h2):(1'h1)] ^ $signed(reg190)) ^ $signed((8'hb1)))} + reg276);
          if ((((^wire196[(2'h3):(1'h1)]) ^ (reg203 ?
              {(reg198 ? (8'hbc) : wire146),
                  (~&reg213)} : $signed(reg251[(4'h8):(2'h3)]))) >= reg263))
            begin
              reg283 <= wire197;
              reg284 <= $signed(wire146[(5'h12):(3'h6)]);
            end
          else
            begin
              reg285 = {(~^reg168[(4'h8):(2'h3)]), reg191[(2'h3):(1'h0)]};
              reg286 <= (~^$signed((reg263[(1'h0):(1'h0)] ?
                  reg187[(1'h1):(1'h0)] : reg233[(3'h7):(3'h6)])));
              reg287 = $unsigned(reg177[(4'hb):(3'h6)]);
            end
        end
      reg288 <= reg276;
      reg289 = ((reg286[(2'h2):(1'h1)] ?
              (({(8'hbe)} && (8'had)) ?
                  ((reg239 == reg234) ?
                      wire149 : $signed(reg212)) : $signed((reg198 ?
                      reg235 : (8'ha4)))) : (((|reg249) ?
                      (reg280 ? reg257 : reg171) : $signed(reg234)) ?
                  ((reg216 ?
                      reg170 : (8'hbd)) >= (reg251 | reg218)) : (8'ha5))) ?
          $signed(reg171) : $unsigned((-(-(reg281 ? reg269 : (8'hb7))))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module30
#(parameter param142 = (~&({(((8'ha9) << (8'haf)) <= (8'hb3)), (!((8'ha1) ? (8'ha4) : (8'hb6)))} <<< (|({(8'hb7), (8'ha8)} != ((8'h9d) ? (8'h9e) : (8'hb2)))))))
(y, clk, wire35, wire34, wire33, wire32, wire31);
  output wire [(32'h50f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire35;
  input wire signed [(4'hf):(1'h0)] wire34;
  input wire [(4'h8):(1'h0)] wire33;
  input wire [(3'h4):(1'h0)] wire32;
  input wire signed [(5'h14):(1'h0)] wire31;
  wire signed [(4'hb):(1'h0)] wire134;
  wire [(5'h10):(1'h0)] wire77;
  wire [(3'h5):(1'h0)] wire76;
  wire signed [(5'h10):(1'h0)] wire75;
  wire [(3'h5):(1'h0)] wire66;
  wire signed [(5'h12):(1'h0)] wire43;
  wire signed [(4'h8):(1'h0)] wire38;
  wire [(5'h12):(1'h0)] wire37;
  wire signed [(5'h14):(1'h0)] wire36;
  reg [(5'h12):(1'h0)] reg141 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg140 = (1'h0);
  reg [(4'hf):(1'h0)] reg139 = (1'h0);
  reg [(4'he):(1'h0)] reg138 = (1'h0);
  reg [(4'hb):(1'h0)] reg137 = (1'h0);
  reg [(3'h6):(1'h0)] reg136 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg135 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg133 = (1'h0);
  reg [(4'ha):(1'h0)] reg131 = (1'h0);
  reg [(4'h9):(1'h0)] reg127 = (1'h0);
  reg [(4'hb):(1'h0)] reg126 = (1'h0);
  reg [(4'h9):(1'h0)] reg125 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg124 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg123 = (1'h0);
  reg [(5'h13):(1'h0)] reg122 = (1'h0);
  reg [(5'h15):(1'h0)] reg121 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg120 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg117 = (1'h0);
  reg [(3'h6):(1'h0)] reg114 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg112 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg110 = (1'h0);
  reg [(2'h2):(1'h0)] reg109 = (1'h0);
  reg [(4'hf):(1'h0)] reg108 = (1'h0);
  reg [(4'ha):(1'h0)] reg107 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg106 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg104 = (1'h0);
  reg [(5'h14):(1'h0)] reg103 = (1'h0);
  reg [(4'hd):(1'h0)] reg101 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg97 = (1'h0);
  reg [(4'hf):(1'h0)] reg100 = (1'h0);
  reg [(4'h9):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg98 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg96 = (1'h0);
  reg [(3'h5):(1'h0)] reg93 = (1'h0);
  reg [(4'h8):(1'h0)] reg92 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg91 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg90 = (1'h0);
  reg signed [(4'he):(1'h0)] reg89 = (1'h0);
  reg [(4'ha):(1'h0)] reg88 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg86 = (1'h0);
  reg [(5'h12):(1'h0)] reg85 = (1'h0);
  reg signed [(4'he):(1'h0)] reg84 = (1'h0);
  reg signed [(4'he):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg82 = (1'h0);
  reg [(3'h7):(1'h0)] reg81 = (1'h0);
  reg [(5'h12):(1'h0)] reg80 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg79 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg74 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg71 = (1'h0);
  reg [(3'h7):(1'h0)] reg70 = (1'h0);
  reg [(5'h12):(1'h0)] reg68 = (1'h0);
  reg [(5'h12):(1'h0)] reg67 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg64 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg63 = (1'h0);
  reg [(4'hb):(1'h0)] reg62 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg57 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg56 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg53 = (1'h0);
  reg [(4'hd):(1'h0)] reg52 = (1'h0);
  reg [(5'h10):(1'h0)] reg51 = (1'h0);
  reg [(5'h11):(1'h0)] reg49 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg48 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg46 = (1'h0);
  reg [(5'h13):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg44 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg42 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg41 = (1'h0);
  reg [(3'h4):(1'h0)] reg40 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg39 = (1'h0);
  reg [(5'h15):(1'h0)] forvar135 = (1'h0);
  reg [(2'h3):(1'h0)] reg132 = (1'h0);
  reg [(4'he):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg129 = (1'h0);
  reg [(5'h14):(1'h0)] reg128 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg119 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar118 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg116 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg115 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar111 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar105 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg102 = (1'h0);
  reg [(4'hf):(1'h0)] forvar97 = (1'h0);
  reg [(4'h9):(1'h0)] reg95 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg94 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg87 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar78 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg73 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg72 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg69 = (1'h0);
  reg [(4'h9):(1'h0)] reg61 = (1'h0);
  reg [(3'h5):(1'h0)] reg60 = (1'h0);
  reg [(2'h3):(1'h0)] reg59 = (1'h0);
  reg [(3'h7):(1'h0)] forvar58 = (1'h0);
  reg [(2'h2):(1'h0)] reg55 = (1'h0);
  reg [(4'h8):(1'h0)] reg54 = (1'h0);
  reg [(4'hb):(1'h0)] forvar51 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg50 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg47 = (1'h0);
  assign y = {wire134,
                 wire77,
                 wire76,
                 wire75,
                 wire66,
                 wire43,
                 wire38,
                 wire37,
                 wire36,
                 reg141,
                 reg140,
                 reg139,
                 reg138,
                 reg137,
                 reg136,
                 reg135,
                 reg133,
                 reg131,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg123,
                 reg122,
                 reg121,
                 reg120,
                 reg117,
                 reg114,
                 reg113,
                 reg112,
                 reg110,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg104,
                 reg103,
                 reg101,
                 reg97,
                 reg100,
                 reg99,
                 reg98,
                 reg96,
                 reg93,
                 reg92,
                 reg91,
                 reg90,
                 reg89,
                 reg88,
                 reg86,
                 reg85,
                 reg84,
                 reg83,
                 reg82,
                 reg81,
                 reg80,
                 reg79,
                 reg74,
                 reg71,
                 reg70,
                 reg68,
                 reg67,
                 reg65,
                 reg64,
                 reg63,
                 reg62,
                 reg57,
                 reg56,
                 reg53,
                 reg52,
                 reg51,
                 reg49,
                 reg48,
                 reg46,
                 reg45,
                 reg44,
                 reg42,
                 reg41,
                 reg40,
                 reg39,
                 forvar135,
                 reg132,
                 reg130,
                 reg129,
                 reg128,
                 reg119,
                 forvar118,
                 reg116,
                 reg115,
                 forvar111,
                 forvar105,
                 reg102,
                 forvar97,
                 reg95,
                 reg94,
                 reg87,
                 forvar78,
                 reg73,
                 reg72,
                 reg69,
                 reg61,
                 reg60,
                 reg59,
                 forvar58,
                 reg55,
                 reg54,
                 forvar51,
                 reg50,
                 reg47,
                 (1'h0)};
  assign wire36 = wire35[(4'he):(3'h6)];
  assign wire37 = wire35[(5'h10):(1'h1)];
  assign wire38 = ($unsigned($signed(wire34)) ?
                      (((!$signed(wire37)) ?
                              (~^(wire31 * wire31)) : ($unsigned(wire35) ^~ ((8'hb5) * (8'hae)))) ?
                          (~&(~(-(8'ha8)))) : $signed($signed($signed(wire31)))) : (&$signed($signed($signed((8'haf))))));
  always
    @(posedge clk) begin
      reg39 <= wire34;
    end
  always
    @(posedge clk) begin
      reg40 <= {$unsigned(((wire34[(4'hf):(4'hd)] || {wire34, wire34}) ?
              wire36[(4'he):(4'h9)] : {(8'haa), wire32[(2'h3):(1'h0)]})),
          (~|($unsigned(wire31[(1'h1):(1'h1)]) < $unsigned((wire37 >> wire33))))};
      reg41 <= ($signed(((wire34 <<< (8'ha3)) ?
              reg39 : $signed((wire33 ? (8'ha1) : wire38)))) ?
          (reg39[(2'h3):(2'h3)] ^ wire34[(3'h6):(3'h6)]) : ($unsigned($unsigned((~|wire34))) && ($signed($signed((8'h9d))) > $unsigned((~reg39)))));
      reg42 <= (((8'h9f) ?
          $signed($unsigned((wire37 & (8'ha2)))) : ((reg40[(2'h2):(2'h2)] ?
                  wire37 : (&reg40)) ?
              $signed((|(8'hb6))) : {(reg41 ?
                      wire36 : wire37)})) + ($signed(reg39[(3'h5):(2'h3)]) | $unsigned($signed((^~reg39)))));
    end
  assign wire43 = $signed(wire33);
  always
    @(posedge clk) begin
      if ((wire32[(2'h3):(1'h0)] <= $signed($unsigned($unsigned($unsigned(wire32))))))
        begin
          reg44 <= (8'ha4);
          reg45 <= wire37;
          reg46 <= ((~^(8'hab)) ?
              (-{wire35[(2'h3):(2'h3)]}) : ((8'hac) ^ wire31[(4'h8):(1'h0)]));
          if ($signed((8'ha1)))
            begin
              reg47 = wire31;
            end
          else
            begin
              reg47 = (8'hb1);
              reg48 <= $unsigned({wire34,
                  (((wire37 - (8'haa)) ? (wire34 | wire31) : (reg47 & wire32)) ?
                      reg41 : reg46)});
            end
        end
      else
        begin
          reg44 <= $unsigned($signed((reg40 + (~^wire32[(2'h2):(1'h0)]))));
          if (((wire32[(1'h1):(1'h1)] ?
              $unsigned($unsigned(reg42[(1'h0):(1'h0)])) : ($signed((wire37 - (8'haf))) && $signed(reg39))) & ((+($unsigned(reg48) ?
              reg47 : (reg45 ?
                  reg40 : wire38))) == ((~&(reg40 != reg39)) < {reg40,
              $signed(reg48)}))))
            begin
              reg45 <= $unsigned(((~|(8'hbb)) ?
                  $unsigned(wire34) : $unsigned($unsigned((~^wire37)))));
              reg46 <= ((reg42 >> $signed($signed((|reg47)))) | $unsigned(wire34[(3'h5):(1'h1)]));
            end
          else
            begin
              reg45 <= wire33[(2'h3):(2'h2)];
            end
          reg48 <= (wire38[(3'h7):(3'h7)] <<< {$unsigned((wire32[(1'h1):(1'h0)] >= {wire36,
                  wire32})),
              $signed($unsigned(wire35[(2'h3):(2'h3)]))});
          if ((wire36 >> (&{($signed(wire36) ~^ {reg45})})))
            begin
              reg49 <= reg42[(3'h6):(1'h0)];
            end
          else
            begin
              reg49 <= $signed(((&($signed(wire34) ?
                      wire38 : (reg49 || wire31))) ?
                  $unsigned($signed(reg42)) : wire37));
            end
          reg50 = wire37;
        end
      if ((8'hbc))
        begin
          reg51 <= wire37[(4'he):(4'he)];
          reg52 <= wire43;
          reg53 <= reg46;
        end
      else
        begin
          for (forvar51 = (1'h0); (forvar51 < (2'h3)); forvar51 = (forvar51 + (1'h1)))
            begin
              reg52 <= (wire33 ?
                  ((($signed(forvar51) ? $signed((8'ha4)) : wire33) ?
                          wire43 : (&{wire37})) ?
                      $unsigned($signed((!wire31))) : ({reg51[(3'h5):(2'h3)]} ?
                          reg44[(1'h0):(1'h0)] : $signed((&wire36)))) : (~^$unsigned(reg50[(1'h1):(1'h0)])));
              reg54 = ($unsigned((~|$signed($signed(wire38)))) >= wire38[(4'h8):(2'h3)]);
              reg55 = $signed({(($unsigned(wire43) & wire38[(3'h7):(3'h5)]) ?
                      ($unsigned(reg49) >>> reg52) : {(reg41 < (8'ha3))})});
            end
          reg56 <= (&reg48);
          reg57 <= reg40[(2'h2):(1'h1)];
          for (forvar58 = (1'h0); (forvar58 < (1'h0)); forvar58 = (forvar58 + (1'h1)))
            begin
              reg59 = wire34[(4'hf):(4'h8)];
              reg60 = ({forvar58,
                      $signed((((7'h40) ?
                          (8'hb3) : wire38) & $signed((8'h9f))))} ?
                  $unsigned($unsigned({(!reg59)})) : (~^wire31));
              reg61 = (reg59 ?
                  reg47[(3'h4):(1'h0)] : {(^$signed((reg48 && reg49)))});
              reg62 <= (((~|reg48) * ($unsigned(reg52[(4'ha):(2'h3)]) ~^ (reg51 && wire31))) ?
                  (reg44 + (|$signed(reg46))) : reg48[(4'ha):(3'h6)]);
              reg63 <= $unsigned((^(((!reg42) && (wire38 != forvar58)) ?
                  $unsigned(reg54) : ((reg60 ? (8'hba) : wire32) ?
                      wire31 : {wire31}))));
            end
          reg64 <= ({forvar51[(1'h0):(1'h0)],
                  $unsigned($signed(wire34[(4'hd):(4'ha)]))} ?
              $unsigned((-reg41[(3'h4):(1'h1)])) : ($signed((&{reg47})) <= reg50[(1'h1):(1'h0)]));
        end
      reg65 <= ({(~(^~reg55))} * forvar51);
    end
  assign wire66 = $unsigned((^~((~&((8'ha8) <= wire32)) ^~ wire31[(3'h4):(2'h3)])));
  always
    @(posedge clk) begin
      if (((&(($signed(wire35) ? reg45 : wire33[(4'h8):(3'h6)]) ?
              reg48[(4'hc):(3'h4)] : (reg42 > $signed(reg65)))) ?
          ((wire35[(4'ha):(1'h1)] ?
              (^(wire32 & reg62)) : $unsigned($unsigned(reg65))) * ($signed($unsigned(reg49)) ^ (((8'h9d) || wire38) && (reg48 + reg65)))) : reg40[(3'h4):(1'h1)]))
        begin
          reg67 <= (~&reg53[(2'h3):(2'h2)]);
          reg68 <= $unsigned($unsigned(reg49[(4'h8):(1'h0)]));
          reg69 = $signed((~&(~&{wire66[(3'h5):(3'h5)]})));
          reg70 <= wire31;
        end
      else
        begin
          reg69 = $signed($unsigned((({reg53, wire38} ?
              (reg39 || reg65) : ((8'hbf) ^~ reg49)) <= (~&wire32))));
        end
    end
  always
    @(posedge clk) begin
      reg71 <= $signed(reg65[(3'h4):(2'h3)]);
      reg72 = {{$signed((~|(wire33 << reg67)))}};
      reg73 = (~$unsigned({$unsigned(reg56)}));
      reg74 <= reg63[(4'he):(3'h7)];
    end
  assign wire75 = ($signed(reg48[(3'h7):(3'h4)]) ~^ $unsigned({$unsigned(reg39[(3'h4):(1'h0)])}));
  assign wire76 = (|{$unsigned(reg57), $unsigned(wire38)});
  assign wire77 = reg74;
  always
    @(posedge clk) begin
      for (forvar78 = (1'h0); (forvar78 < (3'h4)); forvar78 = (forvar78 + (1'h1)))
        begin
          if (((~&reg62) ~^ {(-$signed((reg41 ? reg44 : forvar78)))}))
            begin
              reg79 <= ($signed((8'hbe)) > (reg74 == $unsigned(wire66[(3'h5):(3'h5)])));
              reg80 <= reg70[(2'h2):(2'h2)];
              reg81 <= $signed(((((reg64 ? wire66 : wire35) ?
                  reg56[(4'h8):(1'h0)] : (~^wire77)) ^~ (wire37[(4'hd):(2'h3)] == ((8'hb1) ?
                  reg44 : reg46))) >= (reg52 ?
                  (&reg80) : $unsigned((wire66 ? wire43 : (8'hba))))));
            end
          else
            begin
              reg79 <= $unsigned(wire32[(2'h3):(1'h0)]);
              reg80 <= $unsigned($unsigned($unsigned(((reg45 <= reg57) ?
                  reg44[(5'h10):(2'h3)] : reg40))));
              reg81 <= $unsigned(((|(8'h9f)) <= ((-(reg62 << reg48)) >> $signed((reg45 >>> wire31)))));
              reg82 <= reg46;
              reg83 <= wire76[(2'h2):(2'h2)];
            end
        end
      if ({((-($signed((8'hab)) ?
              wire75[(4'hc):(4'h8)] : $signed(reg67))) >= {(reg48 ?
                  forvar78[(3'h5):(3'h5)] : (-reg39))}),
          reg42[(1'h1):(1'h1)]})
        begin
          reg84 <= reg46[(3'h7):(3'h7)];
          reg85 <= reg40[(1'h1):(1'h0)];
          reg86 <= ({reg52} >>> (~|(&$signed($unsigned(reg48)))));
        end
      else
        begin
          reg84 <= $signed(reg52[(4'hb):(3'h7)]);
          if ((+$signed(reg68[(4'ha):(3'h7)])))
            begin
              reg85 <= (-wire43);
              reg87 = {$signed(($signed($unsigned((8'hae))) ^~ (reg81 <= $signed(wire66))))};
            end
          else
            begin
              reg87 = reg84;
              reg88 <= $unsigned({{((wire76 + reg40) ?
                          (reg57 ~^ reg44) : $unsigned((8'ha8)))},
                  reg63[(4'hb):(2'h2)]});
              reg89 <= (~^(&({forvar78[(3'h6):(1'h1)]} ?
                  ((reg81 >= wire66) - (reg88 - reg49)) : reg64)));
              reg90 <= (!{(-reg52), wire77[(4'he):(2'h2)]});
            end
        end
      reg91 <= (8'hb6);
    end
  always
    @(posedge clk) begin
      reg92 <= $unsigned((+wire43[(4'ha):(1'h1)]));
      reg93 <= $unsigned((-{(((8'hbe) - reg40) ?
              {reg41, (8'hb8)} : reg62[(3'h4):(2'h3)]),
          ((~^reg71) | reg81[(1'h1):(1'h1)])}));
      reg94 = $signed(($signed({(reg62 < reg52)}) ?
          ($unsigned((reg91 ?
              reg44 : reg65)) * reg63[(2'h3):(2'h3)]) : $signed({$unsigned((7'h44))})));
      if ($unsigned((^~(reg93[(3'h4):(1'h0)] ?
          $unsigned(wire37) : $signed(((7'h43) ^ (8'hbf)))))))
        begin
          reg95 = $signed($unsigned((-reg88)));
          reg96 <= {$signed(((8'hae) >= {$signed(wire66), $signed(reg81)})),
              $unsigned(wire76)};
          for (forvar97 = (1'h0); (forvar97 < (2'h2)); forvar97 = (forvar97 + (1'h1)))
            begin
              reg98 <= (^((^~(reg91[(3'h4):(2'h2)] ?
                  $signed(wire76) : (8'ha9))) <= $signed(((reg95 < reg44) > (reg79 ?
                  (8'hab) : reg82)))));
              reg99 <= ((^~(~^(~|(reg82 ? wire66 : wire35)))) >> (-(wire33 ?
                  $signed($signed(wire34)) : ((~^reg48) ?
                      {reg40} : $unsigned(reg65)))));
              reg100 <= ((^~reg71) == ((^{(!reg79), (^reg94)}) && reg64));
            end
        end
      else
        begin
          reg96 <= $signed($signed(({(~&wire35), (~(8'hbc))} > {{reg49},
              reg84[(4'ha):(2'h2)]})));
          reg97 <= reg42;
        end
    end
  always
    @(posedge clk) begin
      reg101 <= ((8'hbd) | $signed($signed($signed(wire36))));
      reg102 = wire31;
      reg103 <= {(&reg86), $signed(reg51)};
      reg104 <= $signed((~|wire31[(4'hb):(3'h7)]));
      for (forvar105 = (1'h0); (forvar105 < (3'h4)); forvar105 = (forvar105 + (1'h1)))
        begin
          if ($signed(($signed($unsigned(reg70[(3'h4):(2'h2)])) >> (~$signed((~|(8'hb3)))))))
            begin
              reg106 <= reg56;
              reg107 <= {reg85};
              reg108 <= reg52[(2'h3):(2'h2)];
              reg109 <= (reg108[(4'h8):(3'h4)] ? wire76 : wire77);
              reg110 <= $signed(((wire37 ?
                  reg44[(4'hc):(3'h5)] : reg48) + ($unsigned(wire31[(4'h8):(3'h4)]) << ($unsigned(reg42) ?
                  {reg82} : $signed(wire32)))));
            end
          else
            begin
              reg106 <= (($signed(((~^reg45) ?
                          (reg41 ? reg104 : (8'ha2)) : reg100)) ?
                      reg82[(4'hc):(1'h1)] : reg45) ?
                  reg108 : {reg106[(4'h8):(4'h8)]});
              reg107 <= reg110;
              reg108 <= $unsigned((~|reg99));
              reg109 <= $signed(reg44[(4'ha):(1'h1)]);
              reg110 <= reg91[(1'h1):(1'h0)];
            end
          for (forvar111 = (1'h0); (forvar111 < (3'h4)); forvar111 = (forvar111 + (1'h1)))
            begin
              reg112 <= ($signed(reg52) ^ ((($unsigned(reg102) ?
                  reg40[(3'h4):(1'h0)] : reg65[(1'h0):(1'h0)]) >= $signed($unsigned(reg96))) || ((wire31 ?
                  $unsigned((8'haa)) : (reg49 <= reg53)) < reg89)));
              reg113 <= ((wire66[(2'h2):(1'h1)] < reg57) >> ($unsigned((~^{(8'ha4)})) <<< $signed((~^{reg103,
                  (7'h42)}))));
              reg114 <= (^~(((|(7'h42)) ?
                  $signed((reg52 ^ wire76)) : ((-reg64) << reg96)) > $signed((7'h40))));
              reg115 = (reg44[(3'h7):(3'h7)] || reg64);
            end
          reg116 = (reg82 ?
              ((((reg114 != wire43) ?
                      (reg45 ? reg52 : reg113) : (reg44 ? forvar105 : wire43)) ?
                  reg85 : reg80[(3'h5):(3'h4)]) <= {{$unsigned(reg109)},
                  reg112}) : reg108);
          reg117 <= wire43[(4'h9):(3'h7)];
        end
    end
  always
    @(posedge clk) begin
      for (forvar118 = (1'h0); (forvar118 < (3'h4)); forvar118 = (forvar118 + (1'h1)))
        begin
          reg119 = $unsigned({reg88, $signed(wire38[(3'h7):(1'h1)])});
          reg120 <= (&reg91[(2'h2):(2'h2)]);
          reg121 <= $signed({(|forvar118)});
          reg122 <= wire38;
          reg123 <= ($signed({(reg63[(1'h0):(1'h0)] ^ {reg103, wire43}),
                  (((8'haa) ? reg70 : wire77) ~^ $unsigned(reg120))}) ?
              $signed(reg79) : (8'hba));
        end
      reg124 <= (8'hb7);
      reg125 <= (~^(wire77[(4'h8):(4'h8)] ? reg67 : wire38[(1'h1):(1'h0)]));
      reg126 <= wire33[(1'h0):(1'h0)];
      if ($unsigned(reg48[(2'h2):(1'h1)]))
        begin
          reg127 <= (~|((($unsigned(reg40) ?
                  (reg63 ? reg100 : reg53) : (~(8'ha5))) <<< $signed({reg88})) ?
              $signed((reg119[(1'h1):(1'h0)] >>> $unsigned(reg67))) : ($unsigned($unsigned(reg64)) ?
                  $signed($unsigned(reg62)) : reg71)));
          if ({(($unsigned((reg53 && (8'haf))) * wire36[(2'h2):(2'h2)]) + ((~|wire66[(3'h4):(2'h3)]) || $signed((8'ha4)))),
              reg57[(4'hb):(3'h7)]})
            begin
              reg128 = (reg46 ?
                  $signed((~((reg97 <= reg126) ?
                      wire76 : $signed(reg121)))) : ((reg124 ?
                          reg117[(4'ha):(2'h3)] : ((|reg93) ?
                              $unsigned(reg53) : $signed(reg83))) ?
                      ((reg113 ? forvar118 : $unsigned((8'haa))) ^ ((reg70 ?
                              (8'h9c) : (8'hb7)) ?
                          (^(8'hb1)) : (8'hb0))) : reg64[(5'h10):(1'h0)]));
              reg129 = (|((-($signed(reg101) ?
                  ((8'hb1) ~^ reg123) : $signed(reg48))) > {(8'ha5), (8'ha6)}));
              reg130 = (+reg57);
            end
          else
            begin
              reg128 = {{(((8'ha9) < (^~reg123)) >>> ((!reg119) ^~ wire77)),
                      ($unsigned(wire34[(4'ha):(2'h2)]) ?
                          $signed($unsigned((8'hb1))) : ({wire66} ?
                              $unsigned((7'h44)) : (wire77 ?
                                  reg57 : (8'ha3))))},
                  reg110[(4'h9):(3'h7)]};
            end
          reg131 <= forvar118[(2'h3):(1'h0)];
          reg132 = reg68;
          reg133 <= ($signed((8'had)) ? reg49[(2'h2):(1'h0)] : (8'haa));
        end
      else
        begin
          reg127 <= wire43;
          reg131 <= $signed($signed($signed($signed($unsigned(wire32)))));
        end
    end
  assign wire134 = ((((!reg49) ?
                           $signed(reg83) : {$signed(wire34)}) << $unsigned({(reg63 ?
                               reg122 : (8'ha9))})) ?
                       reg107[(4'h8):(2'h3)] : ({reg80[(3'h6):(3'h4)],
                               reg85[(3'h6):(2'h3)]} ?
                           (reg100[(4'hc):(1'h0)] != ((reg64 ?
                                   wire66 : (8'hb3)) ?
                               (^(7'h40)) : $signed(reg104))) : {{reg62[(4'hb):(2'h3)],
                                   reg82[(4'hd):(2'h2)]},
                               {reg133, ((8'ha4) ? reg40 : reg81)}}));
  always
    @(posedge clk) begin
      if ((^~reg68[(4'hb):(2'h3)]))
        begin
          reg135 <= (&reg83[(1'h0):(1'h0)]);
        end
      else
        begin
          for (forvar135 = (1'h0); (forvar135 < (1'h1)); forvar135 = (forvar135 + (1'h1)))
            begin
              reg136 <= ($signed(reg99[(1'h0):(1'h0)]) << $signed(($unsigned(reg57[(1'h0):(1'h0)]) ?
                  (-((8'h9d) ? wire36 : reg64)) : (reg48 - (reg124 ?
                      reg125 : wire38)))));
              reg137 <= ($unsigned(($signed($unsigned(reg121)) ?
                      reg41 : $unsigned($unsigned(wire34)))) ?
                  wire36 : $signed({wire76[(2'h3):(2'h2)]}));
              reg138 <= (reg97 * $signed((reg57[(5'h10):(4'h8)] + reg88)));
              reg139 <= reg63[(4'hb):(3'h7)];
            end
          reg140 <= (^(((^~(wire76 <<< reg65)) >= $unsigned($unsigned(reg83))) ?
              reg86 : reg81[(2'h3):(1'h0)]));
          reg141 <= (+reg106[(5'h13):(1'h0)]);
        end
    end
endmodule