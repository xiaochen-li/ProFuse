(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h1d9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h2):(1'h0)] wire0;
  input wire signed [(5'h13):(1'h0)] wire1;
  input wire signed [(5'h10):(1'h0)] wire2;
  input wire signed [(4'hd):(1'h0)] wire3;
  wire signed [(5'h13):(1'h0)] wire269;
  wire [(5'h12):(1'h0)] wire268;
  wire signed [(5'h14):(1'h0)] wire267;
  wire [(3'h4):(1'h0)] wire33;
  wire [(4'h8):(1'h0)] wire39;
  wire [(5'h10):(1'h0)] wire40;
  wire [(3'h5):(1'h0)] wire41;
  wire signed [(4'hc):(1'h0)] wire116;
  wire signed [(5'h14):(1'h0)] wire131;
  wire signed [(3'h4):(1'h0)] wire265;
  reg signed [(4'he):(1'h0)] reg128 = (1'h0);
  reg [(4'hc):(1'h0)] reg127 = (1'h0);
  reg [(3'h6):(1'h0)] reg126 = (1'h0);
  reg [(4'he):(1'h0)] reg125 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg124 = (1'h0);
  reg [(4'he):(1'h0)] reg121 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg118 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg38 = (1'h0);
  reg [(5'h11):(1'h0)] reg36 = (1'h0);
  reg [(3'h7):(1'h0)] reg35 = (1'h0);
  reg [(5'h14):(1'h0)] reg14 = (1'h0);
  reg [(5'h10):(1'h0)] reg13 = (1'h0);
  reg [(5'h15):(1'h0)] reg12 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg11 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg10 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg8 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg7 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg6 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg130 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar129 = (1'h0);
  reg signed [(4'he):(1'h0)] reg123 = (1'h0);
  reg [(5'h12):(1'h0)] forvar122 = (1'h0);
  reg [(2'h3):(1'h0)] forvar120 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar119 = (1'h0);
  reg [(5'h11):(1'h0)] reg37 = (1'h0);
  reg [(5'h12):(1'h0)] forvar9 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar5 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar4 = (1'h0);
  assign y = {wire269,
                 wire268,
                 wire267,
                 wire33,
                 wire39,
                 wire40,
                 wire41,
                 wire116,
                 wire131,
                 wire265,
                 reg128,
                 reg127,
                 reg126,
                 reg125,
                 reg124,
                 reg121,
                 reg118,
                 reg38,
                 reg36,
                 reg35,
                 reg14,
                 reg13,
                 reg12,
                 reg11,
                 reg10,
                 reg8,
                 reg7,
                 reg6,
                 reg130,
                 forvar129,
                 reg123,
                 forvar122,
                 forvar120,
                 forvar119,
                 reg37,
                 forvar9,
                 forvar5,
                 forvar4,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar4 = (1'h0); (forvar4 < (3'h4)); forvar4 = (forvar4 + (1'h1)))
        begin
          for (forvar5 = (1'h0); (forvar5 < (2'h3)); forvar5 = (forvar5 + (1'h1)))
            begin
              reg6 <= (8'ha5);
            end
          reg7 <= $unsigned((wire3 ?
              wire1[(3'h7):(3'h7)] : wire2[(4'hd):(4'hc)]));
          reg8 <= $signed((reg6 >>> $unsigned(reg7[(2'h2):(1'h0)])));
          for (forvar9 = (1'h0); (forvar9 < (2'h2)); forvar9 = (forvar9 + (1'h1)))
            begin
              reg10 <= wire2[(3'h6):(2'h3)];
              reg11 <= reg8;
              reg12 <= wire0;
            end
        end
      reg13 <= (8'hbc);
      reg14 <= wire3[(2'h3):(1'h1)];
    end
  module15 #() modinst34 (.wire17(wire1), .clk(clk), .wire16(wire2), .wire19(reg14), .wire18(reg13), .y(wire33));
  always
    @(posedge clk) begin
      reg35 <= $unsigned(($unsigned(reg12[(4'hd):(4'hb)]) & wire3));
      reg36 <= $unsigned(reg14[(1'h0):(1'h0)]);
      reg37 = reg36;
      reg38 <= (+$signed(reg6[(3'h7):(2'h2)]));
    end
  assign wire39 = $signed(reg36);
  assign wire40 = reg12;
  assign wire41 = $unsigned(($signed($unsigned(((8'hb9) ?
                      (7'h41) : wire39))) & reg14[(4'ha):(1'h0)]));
  module42 #() modinst117 (wire116, clk, reg14, reg36, wire40, wire3);
  always
    @(posedge clk) begin
      reg118 <= wire3[(2'h2):(1'h0)];
      for (forvar119 = (1'h0); (forvar119 < (3'h4)); forvar119 = (forvar119 + (1'h1)))
        begin
          for (forvar120 = (1'h0); (forvar120 < (1'h0)); forvar120 = (forvar120 + (1'h1)))
            begin
              reg121 <= ((wire0[(1'h0):(1'h0)] ?
                  {$unsigned({reg10,
                          wire3})} : (-((^forvar119) ^ (wire39 <= wire33)))) ~^ (~&$unsigned(reg10)));
            end
          for (forvar122 = (1'h0); (forvar122 < (1'h0)); forvar122 = (forvar122 + (1'h1)))
            begin
              reg123 = wire1;
            end
          reg124 <= forvar122[(4'hb):(3'h6)];
          reg125 <= $unsigned((+(reg7[(3'h4):(2'h3)] ?
              $signed((reg35 ? wire116 : reg12)) : forvar120[(2'h3):(2'h3)])));
          reg126 <= $unsigned((!reg124));
        end
      reg127 <= $unsigned((&({$signed(forvar122), (^(8'haa))} ?
          $signed((wire3 ? (7'h43) : reg6)) : (reg11 ?
              $unsigned((8'h9f)) : wire3[(3'h4):(3'h4)]))));
      reg128 <= $unsigned(((~^$unsigned(reg14[(5'h10):(1'h1)])) ?
          $unsigned($unsigned($signed((8'haa)))) : (-$signed((8'hb2)))));
      for (forvar129 = (1'h0); (forvar129 < (1'h0)); forvar129 = (forvar129 + (1'h1)))
        begin
          reg130 = $unsigned({reg12[(1'h1):(1'h0)]});
        end
    end
  assign wire131 = {reg14[(5'h10):(4'he)],
                       ((^reg124[(2'h2):(2'h2)]) >= wire116[(1'h0):(1'h0)])};
  module132 #() modinst266 (wire265, clk, reg12, reg127, reg126, reg13, wire116);
  assign wire267 = $unsigned(((+$unsigned($signed((8'hbf)))) ?
                       $signed({((8'hb8) + reg118),
                           wire40[(4'h8):(4'h8)]}) : $unsigned($signed($unsigned(reg10)))));
  assign wire268 = ((~($signed($unsigned(wire267)) ?
                       $unsigned($signed((8'hab))) : $unsigned((reg6 >= wire265)))) <= ($signed((wire267 ?
                       wire265 : $signed(reg10))) | (~|($unsigned(wire265) != reg8))));
  assign wire269 = reg126[(2'h3):(2'h2)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module132
#(parameter param264 = (((8'h9e) ? (^{((8'hbe) << (8'hb7))}) : (+(((8'ha2) == (8'ha8)) ? (8'hb6) : (~|(8'haa))))) ? (8'hac) : ((^(^{(8'hb9)})) ? (-(~^{(8'h9c)})) : (~|{((8'hb0) >> (8'ha8)), ((8'hbf) ? (7'h44) : (8'hb6))}))))
(y, clk, wire137, wire136, wire135, wire134, wire133);
  output wire [(32'h22c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'he):(1'h0)] wire137;
  input wire [(4'hc):(1'h0)] wire136;
  input wire [(3'h6):(1'h0)] wire135;
  input wire signed [(4'he):(1'h0)] wire134;
  input wire [(4'hc):(1'h0)] wire133;
  wire signed [(4'h8):(1'h0)] wire263;
  wire signed [(4'he):(1'h0)] wire262;
  wire signed [(2'h3):(1'h0)] wire260;
  wire signed [(3'h4):(1'h0)] wire245;
  wire signed [(3'h6):(1'h0)] wire244;
  wire signed [(4'hf):(1'h0)] wire184;
  wire [(5'h12):(1'h0)] wire172;
  wire [(3'h7):(1'h0)] wire142;
  wire signed [(4'h8):(1'h0)] wire138;
  wire signed [(4'he):(1'h0)] wire242;
  reg signed [(5'h12):(1'h0)] reg171 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg170 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg169 = (1'h0);
  reg [(5'h12):(1'h0)] reg168 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg167 = (1'h0);
  reg signed [(4'he):(1'h0)] reg166 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg163 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg159 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg161 = (1'h0);
  reg signed [(4'he):(1'h0)] reg160 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg158 = (1'h0);
  reg [(4'h9):(1'h0)] reg157 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg156 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg153 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg152 = (1'h0);
  reg [(3'h5):(1'h0)] reg151 = (1'h0);
  reg [(5'h14):(1'h0)] reg150 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg149 = (1'h0);
  reg [(4'he):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg147 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg145 = (1'h0);
  reg signed [(4'he):(1'h0)] reg144 = (1'h0);
  reg [(4'he):(1'h0)] reg143 = (1'h0);
  reg [(5'h10):(1'h0)] reg141 = (1'h0);
  reg [(5'h14):(1'h0)] reg140 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg139 = (1'h0);
  reg [(3'h4):(1'h0)] reg165 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar160 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg162 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar159 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg155 = (1'h0);
  reg [(5'h10):(1'h0)] forvar154 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg146 = (1'h0);
  assign y = {wire263,
                 wire262,
                 wire260,
                 wire245,
                 wire244,
                 wire184,
                 wire172,
                 wire142,
                 wire138,
                 wire242,
                 reg171,
                 reg170,
                 reg169,
                 reg168,
                 reg167,
                 reg166,
                 reg164,
                 reg163,
                 reg159,
                 reg161,
                 reg160,
                 reg158,
                 reg157,
                 reg156,
                 reg153,
                 reg152,
                 reg151,
                 reg150,
                 reg149,
                 reg148,
                 reg147,
                 reg145,
                 reg144,
                 reg143,
                 reg141,
                 reg140,
                 reg139,
                 reg165,
                 forvar160,
                 reg162,
                 forvar159,
                 reg155,
                 forvar154,
                 reg146,
                 (1'h0)};
  assign wire138 = (^wire135[(3'h6):(2'h3)]);
  always
    @(posedge clk) begin
      reg139 <= $unsigned((wire133[(4'h8):(2'h2)] ?
          wire133[(4'h9):(4'h8)] : $unsigned($signed((wire137 ?
              wire138 : wire134)))));
      reg140 <= wire135[(3'h6):(3'h6)];
      reg141 <= (^$signed((~{reg139[(1'h0):(1'h0)], reg139[(3'h5):(3'h5)]})));
    end
  assign wire142 = wire138;
  always
    @(posedge clk) begin
      reg143 <= {($signed($unsigned((wire137 ? reg140 : reg140))) ?
              ($unsigned((wire133 | wire137)) ?
                  wire136[(2'h2):(2'h2)] : $signed((wire138 && (8'hb7)))) : wire133),
          wire134};
      if (reg139[(1'h0):(1'h0)])
        begin
          if ($unsigned(($unsigned(wire137) ~^ {$unsigned((wire137 > reg143))})))
            begin
              reg144 <= $signed((|((|reg139[(1'h1):(1'h1)]) & $signed((|(8'hab))))));
            end
          else
            begin
              reg144 <= (^~(8'ha5));
              reg145 <= $unsigned($signed((!{(reg144 < wire137),
                  $unsigned(wire137)})));
              reg146 = wire138;
              reg147 <= (({($unsigned(wire133) * {reg139})} ?
                  reg145[(5'h12):(4'hd)] : ((reg145[(4'h8):(4'h8)] + reg144) ?
                      $unsigned(wire137) : $unsigned({wire137,
                          (8'haf)}))) != $unsigned((($signed(reg141) ?
                  (&wire136) : $signed(wire138)) == (reg139[(2'h3):(1'h0)] ?
                  reg141[(2'h2):(2'h2)] : $signed(reg145)))));
              reg148 <= $signed(($unsigned((reg144 ?
                  reg141 : reg141)) > reg147));
            end
          reg149 <= ($signed((wire142[(2'h3):(1'h1)] ?
                  (^~wire133[(3'h4):(1'h0)]) : wire133[(3'h6):(2'h2)])) ?
              (reg145[(3'h7):(3'h5)] ?
                  $unsigned(reg146[(1'h1):(1'h0)]) : wire138[(2'h2):(2'h2)]) : $signed(reg146));
        end
      else
        begin
          if ({(reg139[(3'h5):(1'h0)] <<< reg141)})
            begin
              reg144 <= (~^$signed($unsigned((8'hbc))));
              reg145 <= ((reg143 ?
                  $signed(((reg149 | reg147) < wire136)) : (|$signed($unsigned(reg148)))) > (((reg139[(4'h8):(1'h0)] ?
                      $unsigned(wire136) : wire135) ?
                  ((-reg148) ? {wire135} : (-wire136)) : (reg144 ?
                      reg148 : (wire135 ?
                          reg149 : reg148))) <<< $signed(((!reg144) < (reg143 ?
                  wire137 : reg145)))));
              reg147 <= reg139;
              reg148 <= reg147;
              reg149 <= reg147[(1'h0):(1'h0)];
            end
          else
            begin
              reg146 = reg145;
              reg147 <= ($unsigned({((wire136 * (8'ha9)) ?
                          $signed(wire134) : (wire135 <= wire133))}) ?
                  reg139 : wire142[(3'h6):(2'h2)]);
            end
          reg150 <= {reg140[(3'h4):(1'h1)], reg139};
          reg151 <= $signed(wire133);
          reg152 <= ($signed({((+wire137) - reg140[(3'h4):(1'h1)]), wire134}) ?
              $signed((^~(((8'hb6) << reg148) ?
                  $unsigned((8'ha0)) : reg140))) : (8'haa));
          reg153 <= (wire134[(1'h1):(1'h0)] - $unsigned({wire134}));
        end
      for (forvar154 = (1'h0); (forvar154 < (2'h3)); forvar154 = (forvar154 + (1'h1)))
        begin
          if ((reg145[(4'hf):(4'h9)] << (((~|reg145[(4'h8):(2'h2)]) ?
              wire138 : reg153) << reg146)))
            begin
              reg155 = {(|$unsigned(wire138))};
            end
          else
            begin
              reg156 <= (~|{$signed($signed({reg140, reg140}))});
              reg157 <= ((+{reg151}) == ({$unsigned(reg153), (~|reg145)} ?
                  $unsigned((^(reg141 ?
                      wire133 : reg152))) : (reg141[(1'h1):(1'h0)] ?
                      wire134[(4'h9):(3'h5)] : $unsigned(reg148))));
            end
        end
      reg158 <= ($signed(((reg149[(2'h3):(1'h1)] ?
          (reg149 ? reg147 : (8'hb3)) : (forvar154 > reg155)) << ((reg139 ?
              reg152 : wire137) ?
          {(8'hae)} : (reg143 ^~ reg149)))) <<< {((wire135 | (~wire135)) ?
              reg157[(1'h1):(1'h1)] : reg149)});
      if (($unsigned(((((8'h9f) ? reg140 : (7'h40)) ?
              (reg158 ? (8'hb0) : reg155) : (reg144 && reg145)) ?
          $signed((reg158 ?
              wire133 : reg152)) : $unsigned(reg149[(4'hf):(4'hd)]))) && reg156))
        begin
          for (forvar159 = (1'h0); (forvar159 < (1'h1)); forvar159 = (forvar159 + (1'h1)))
            begin
              reg160 <= (!forvar154[(4'hd):(4'hd)]);
              reg161 <= {(&(+$signed($unsigned(reg158))))};
              reg162 = ((reg155 ?
                  reg139 : reg156[(1'h0):(1'h0)]) & (forvar154[(4'he):(4'ha)] || wire136[(4'hb):(3'h5)]));
            end
        end
      else
        begin
          reg159 <= (reg141 * (((&((8'hb6) == wire134)) >>> ({(8'hae), reg147} ?
                  forvar159[(4'he):(3'h5)] : forvar159)) ?
              (-(^~(|forvar154))) : (^~$signed((7'h42)))));
          for (forvar160 = (1'h0); (forvar160 < (3'h4)); forvar160 = (forvar160 + (1'h1)))
            begin
              reg162 = reg141[(2'h2):(1'h0)];
              reg163 <= $unsigned(wire135[(1'h0):(1'h0)]);
              reg164 <= (({{((7'h41) ?
                          reg159 : forvar154)}} ^~ wire137) == (7'h41));
              reg165 = reg140[(4'h8):(1'h1)];
            end
          reg166 <= ((~|(reg157 <= wire134[(4'h9):(3'h7)])) ?
              reg160 : ((~|reg143) ?
                  $signed(wire133[(2'h2):(1'h1)]) : $unsigned($signed((reg158 ?
                      wire135 : reg161)))));
          reg167 <= reg147[(1'h0):(1'h0)];
          if ((!reg150[(4'hf):(1'h1)]))
            begin
              reg168 <= reg159;
              reg169 <= wire134[(2'h3):(1'h0)];
              reg170 <= ((^(((~^(8'hb4)) || reg167[(2'h2):(1'h1)]) ?
                      reg162 : $unsigned(reg162[(3'h6):(3'h6)]))) ?
                  ($signed($signed(((8'h9e) ?
                      reg146 : reg162))) ^~ (reg155[(3'h7):(3'h4)] < ($unsigned(forvar159) ?
                      $unsigned(reg147) : $signed(reg149)))) : (reg160 <<< (reg165[(3'h4):(1'h0)] & $unsigned((wire137 ?
                      wire135 : wire137)))));
              reg171 <= reg141[(3'h5):(2'h2)];
            end
          else
            begin
              reg168 <= $unsigned(reg167);
              reg169 <= reg147;
            end
        end
    end
  assign wire172 = reg153[(1'h1):(1'h1)];
  module173 #() modinst185 (wire184, clk, wire142, reg140, reg157, reg152, reg158);
  module186 #() modinst243 (.y(wire242), .wire187(reg159), .wire189(reg160), .clk(clk), .wire190(wire134), .wire188(reg171));
  assign wire244 = ($unsigned((((wire133 * reg168) < {reg144,
                       reg143}) >= ($signed(wire184) ?
                       reg163[(1'h0):(1'h0)] : $signed(wire184)))) ^ (~|reg140[(1'h0):(1'h0)]));
  assign wire245 = ((^~$unsigned(reg170)) == $signed($signed(reg170)));
  module246 #() modinst261 (wire260, clk, reg152, reg141, reg147, reg160, reg139);
  assign wire262 = (-{(!wire242[(2'h2):(1'h1)])});
  assign wire263 = wire136[(3'h7):(1'h0)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module42
#(parameter param115 = ((((((7'h41) ? (8'hbb) : (7'h41)) < ((8'ha6) < (8'haa))) ? (!((8'ha9) ? (8'hb6) : (8'hb1))) : {(^(8'h9d))}) ^~ (^(((8'ha5) != (8'hab)) ? (+(8'ha2)) : ((8'hae) ? (8'h9c) : (7'h44))))) ~^ (({(~&(8'hb1)), {(8'hbf)}} <= ((~^(8'hbf)) >= ((8'had) ? (8'hab) : (8'hac)))) ~^ ({((8'hae) ? (8'hb8) : (8'hb3)), {(8'hb1), (8'hba)}} ? (~|((7'h42) <= (8'ha6))) : ({(8'hab), (8'ha9)} ? ((8'hae) << (8'ha9)) : ((8'h9c) == (8'hbd)))))))
(y, clk, wire46, wire45, wire44, wire43);
  output wire [(32'h78):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h14):(1'h0)] wire46;
  input wire [(5'h11):(1'h0)] wire45;
  input wire [(5'h10):(1'h0)] wire44;
  input wire signed [(4'hd):(1'h0)] wire43;
  wire signed [(4'he):(1'h0)] wire114;
  wire signed [(5'h11):(1'h0)] wire113;
  wire signed [(5'h13):(1'h0)] wire112;
  wire signed [(5'h12):(1'h0)] wire77;
  wire signed [(5'h14):(1'h0)] wire48;
  wire signed [(5'h12):(1'h0)] wire47;
  wire [(4'hd):(1'h0)] wire110;
  assign y = {wire114,
                 wire113,
                 wire112,
                 wire77,
                 wire48,
                 wire47,
                 wire110,
                 (1'h0)};
  assign wire47 = (wire44 ?
                      wire43[(4'h8):(2'h3)] : ((~|wire45[(4'hc):(3'h7)]) != wire45));
  assign wire48 = wire44[(1'h1):(1'h0)];
  module49 #() modinst78 (.wire52(wire45), .wire53(wire43), .clk(clk), .wire50(wire47), .y(wire77), .wire51(wire46), .wire54(wire44));
  module79 #() modinst111 (.wire80(wire45), .y(wire110), .wire81(wire77), .clk(clk), .wire82(wire43), .wire84(wire48), .wire83(wire44));
  assign wire112 = (!(($unsigned(wire45[(4'hc):(4'ha)]) ?
                           ({wire47} ?
                               (wire47 >>> wire48) : $signed(wire48)) : wire43[(2'h2):(1'h0)]) ?
                       (((~(8'hb2)) ?
                               (wire46 ?
                                   wire48 : wire44) : wire44[(4'he):(2'h3)]) ?
                           {$signed(wire77)} : $signed(wire44[(4'hb):(2'h3)])) : (($signed(wire43) ?
                               (wire43 ? (8'hb8) : wire77) : (wire43 ?
                                   wire47 : (8'ha5))) ?
                           (wire77[(4'hf):(4'he)] | wire45) : ({wire77,
                               wire46} <= wire48[(4'h9):(4'h9)]))));
  assign wire113 = wire48;
  assign wire114 = {((&$unsigned((~|wire112))) ?
                           $unsigned({wire45,
                               ((8'hb5) == wire46)}) : $signed((!wire46[(5'h13):(1'h0)]))),
                       $signed(($unsigned((wire47 << (8'ha9))) ?
                           (wire47[(3'h7):(1'h1)] - (+(8'hab))) : wire47))};
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module15  (y, clk, wire19, wire18, wire17, wire16);
  output wire [(32'h8c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h11):(1'h0)] wire19;
  input wire signed [(3'h7):(1'h0)] wire18;
  input wire signed [(5'h13):(1'h0)] wire17;
  input wire [(4'hb):(1'h0)] wire16;
  wire [(5'h12):(1'h0)] wire21;
  wire [(3'h5):(1'h0)] wire20;
  reg [(4'he):(1'h0)] reg31 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg30 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg23 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg28 = (1'h0);
  reg [(5'h10):(1'h0)] reg27 = (1'h0);
  reg [(3'h5):(1'h0)] reg26 = (1'h0);
  reg [(3'h6):(1'h0)] reg25 = (1'h0);
  reg [(3'h7):(1'h0)] reg24 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg32 = (1'h0);
  reg [(2'h2):(1'h0)] reg29 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar22 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar23 = (1'h0);
  reg [(3'h6):(1'h0)] reg22 = (1'h0);
  assign y = {wire21,
                 wire20,
                 reg31,
                 reg30,
                 reg23,
                 reg28,
                 reg27,
                 reg26,
                 reg25,
                 reg24,
                 reg32,
                 reg29,
                 forvar22,
                 forvar23,
                 reg22,
                 (1'h0)};
  assign wire20 = wire19;
  assign wire21 = $unsigned($unsigned(wire17[(1'h1):(1'h0)]));
  always
    @(posedge clk) begin
      if ({$signed(wire19), wire17})
        begin
          reg22 = wire21[(4'hd):(3'h5)];
          for (forvar23 = (1'h0); (forvar23 < (1'h1)); forvar23 = (forvar23 + (1'h1)))
            begin
              reg24 <= wire17;
              reg25 <= reg22[(2'h2):(1'h1)];
              reg26 <= wire19;
              reg27 <= ($signed(((wire20[(1'h1):(1'h0)] <<< {wire17}) & forvar23[(3'h7):(3'h6)])) << (~^({(-wire17),
                  $signed(wire18)} * wire21[(1'h1):(1'h0)])));
            end
          reg28 <= $signed((($unsigned(forvar23) <<< (|reg27[(4'hc):(3'h6)])) ~^ (reg25[(1'h0):(1'h0)] ?
              (reg24[(2'h3):(1'h1)] ?
                  (8'h9d) : $unsigned(wire17)) : wire19[(4'hc):(4'h8)])));
        end
      else
        begin
          for (forvar22 = (1'h0); (forvar22 < (3'h4)); forvar22 = (forvar22 + (1'h1)))
            begin
              reg23 <= ($unsigned($unsigned(($unsigned(reg22) ?
                  (wire18 != wire16) : (wire20 <= reg26)))) == $unsigned((^~(8'ha4))));
              reg24 <= wire16[(3'h4):(3'h4)];
              reg29 = $unsigned(reg26);
              reg30 <= (reg25[(2'h2):(2'h2)] != (^wire18[(2'h3):(1'h1)]));
              reg31 <= $unsigned($signed($unsigned(($signed(reg28) > {(8'haa)}))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg32 = ($signed(wire20[(2'h3):(2'h3)]) >>> (((reg27[(5'h10):(4'ha)] >>> {reg25,
              reg28}) && ($signed(reg30) ~^ (reg23 ? (8'hb6) : wire20))) ?
          ((+{wire20, wire16}) ?
              (!(wire21 ? reg25 : (8'hbd))) : ((&reg31) ?
                  (^~wire19) : (wire21 ?
                      reg26 : wire19))) : $signed({(~|reg30)})));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module79
#(parameter param108 = {(({((8'hbb) ? (7'h43) : (8'hb1)), {(8'hb5), (8'hb0)}} ? (((7'h44) ? (7'h40) : (8'h9e)) ? ((8'h9d) | (8'h9d)) : (8'hac)) : (((8'hb6) ~^ (8'hb9)) ? ((7'h42) - (8'haa)) : (^(8'hbe)))) ? ((((8'haf) ? (8'hba) : (8'hb7)) ? (~|(8'hbc)) : ((8'hb5) || (7'h41))) ? (|((8'hb3) ? (8'hab) : (8'ha8))) : {((8'ha4) == (8'hb7)), ((8'hb1) ? (8'hb3) : (8'h9f))}) : ((((8'had) - (8'ha0)) > {(8'ha7)}) >= (8'hbc)))}, 
parameter param109 = {(param108 ? param108 : (param108 ? param108 : param108))})
(y, clk, wire84, wire83, wire82, wire81, wire80);
  output wire [(32'heb):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h14):(1'h0)] wire84;
  input wire [(3'h7):(1'h0)] wire83;
  input wire [(4'hd):(1'h0)] wire82;
  input wire signed [(3'h7):(1'h0)] wire81;
  input wire [(3'h6):(1'h0)] wire80;
  wire signed [(2'h2):(1'h0)] wire90;
  wire signed [(5'h12):(1'h0)] wire89;
  wire signed [(5'h15):(1'h0)] wire88;
  wire signed [(2'h2):(1'h0)] wire86;
  wire [(3'h5):(1'h0)] wire85;
  reg [(4'h9):(1'h0)] reg107 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg106 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg103 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg102 = (1'h0);
  reg [(3'h6):(1'h0)] reg99 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg96 = (1'h0);
  reg [(4'hb):(1'h0)] reg95 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg93 = (1'h0);
  reg [(2'h3):(1'h0)] reg92 = (1'h0);
  reg [(4'h8):(1'h0)] reg91 = (1'h0);
  reg [(4'he):(1'h0)] reg105 = (1'h0);
  reg [(5'h13):(1'h0)] reg104 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg101 = (1'h0);
  reg [(2'h2):(1'h0)] reg100 = (1'h0);
  reg [(4'h8):(1'h0)] forvar98 = (1'h0);
  reg [(5'h13):(1'h0)] reg97 = (1'h0);
  reg [(4'h9):(1'h0)] reg94 = (1'h0);
  reg [(4'hf):(1'h0)] forvar94 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg87 = (1'h0);
  assign y = {wire90,
                 wire89,
                 wire88,
                 wire86,
                 wire85,
                 reg107,
                 reg106,
                 reg103,
                 reg102,
                 reg99,
                 reg96,
                 reg95,
                 reg93,
                 reg92,
                 reg91,
                 reg105,
                 reg104,
                 reg101,
                 reg100,
                 forvar98,
                 reg97,
                 reg94,
                 forvar94,
                 reg87,
                 (1'h0)};
  assign wire85 = wire80[(3'h5):(1'h0)];
  assign wire86 = wire81;
  always
    @(posedge clk) begin
      reg87 = {(8'hbd)};
    end
  assign wire88 = $signed((+wire80));
  assign wire89 = (-(($unsigned(wire81[(3'h5):(3'h4)]) ?
                          ($signed(wire83) >= {wire86}) : ((&wire80) + (wire84 <<< wire86))) ?
                      {(^~$signed(wire82)),
                          (wire81[(3'h4):(1'h1)] ?
                              (wire82 ?
                                  wire80 : wire85) : (&(8'hbd)))} : (((wire84 <<< wire82) ?
                              wire86[(1'h1):(1'h1)] : (wire80 | (8'ha9))) ?
                          $unsigned((wire86 >>> wire85)) : wire81)));
  assign wire90 = {$unsigned({($signed(wire85) == {wire89})})};
  always
    @(posedge clk) begin
      reg91 <= $unsigned((8'hb7));
      reg92 <= wire85;
    end
  always
    @(posedge clk) begin
      if ($signed(({$signed((wire81 <<< wire85)), (^~$unsigned((8'ha5)))} ?
          (-$unsigned((wire81 ?
              wire85 : (7'h44)))) : ((+(wire85 >>> reg91)) ^ wire84))))
        begin
          reg93 <= {$signed($unsigned(((wire89 & wire83) < wire83[(2'h2):(1'h0)]))),
              wire81[(3'h5):(3'h4)]};
          for (forvar94 = (1'h0); (forvar94 < (2'h3)); forvar94 = (forvar94 + (1'h1)))
            begin
              reg95 <= $unsigned(($unsigned((+$unsigned(reg92))) ?
                  $unsigned($signed((!wire82))) : (-(|((8'hb8) - wire85)))));
            end
          reg96 <= ((~reg91) == wire80[(3'h4):(2'h3)]);
        end
      else
        begin
          reg93 <= (-$unsigned(({((8'ha3) ? (8'ha9) : reg95)} ?
              (8'hbe) : ((reg96 * wire81) << $signed(wire83)))));
          if (((~$unsigned(($signed(forvar94) ?
                  $signed(forvar94) : (reg95 + wire81)))) ?
              ((reg92 >= forvar94) ?
                  ($signed($signed(reg92)) ?
                      ((wire86 | reg96) ~^ (~&wire81)) : (forvar94 >>> {forvar94,
                          wire81})) : wire83[(3'h4):(1'h0)]) : {$signed(((~&wire81) >= $signed(wire81))),
                  (^~wire88[(3'h7):(3'h6)])}))
            begin
              reg94 = (reg96[(4'h8):(3'h5)] >> reg96);
            end
          else
            begin
              reg94 = $unsigned($signed($signed({$unsigned((7'h43))})));
            end
          reg95 <= wire88;
          reg97 = {wire82[(4'h9):(4'h8)],
              (({((8'ha0) ? wire89 : wire81)} ?
                      wire85 : (((8'h9f) ?
                          wire82 : wire82) == forvar94[(3'h4):(1'h0)])) ?
                  $unsigned(((reg94 || forvar94) ?
                      $signed(reg96) : (wire90 ?
                          wire88 : reg92))) : ($unsigned((8'ha9)) ?
                      $signed(wire89) : (wire82 > ((8'ha6) >> reg92))))};
          for (forvar98 = (1'h0); (forvar98 < (2'h3)); forvar98 = (forvar98 + (1'h1)))
            begin
              reg99 <= ((^~reg96) ?
                  ({$unsigned((reg97 ? reg95 : reg94))} ?
                      (wire88 ?
                          $signed({(7'h43),
                              reg97}) : ((~&wire80) ~^ (^forvar94))) : wire83[(2'h3):(1'h0)]) : wire84[(2'h3):(2'h3)]);
              reg100 = wire85[(1'h0):(1'h0)];
              reg101 = $unsigned(wire83[(2'h3):(1'h0)]);
              reg102 <= $unsigned($unsigned(($unsigned((-wire80)) ?
                  (8'hb7) : {$unsigned((7'h44))})));
              reg103 <= $signed(((^~wire83) ? forvar94 : reg97[(1'h0):(1'h0)]));
            end
        end
      reg104 = reg97[(4'hd):(3'h4)];
      reg105 = $signed($signed(wire89[(5'h10):(4'he)]));
      reg106 <= $signed($signed(reg101[(3'h6):(1'h0)]));
      reg107 <= (^$signed(($signed(wire88) ?
          $signed((reg101 ^ reg94)) : reg93)));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module49
#(parameter param76 = (({({(7'h43), (8'hbe)} ? (~&(8'h9f)) : (8'hac)), (~&((7'h41) != (7'h43)))} - (((-(8'hb3)) ? {(7'h43), (8'ha1)} : ((8'ha7) ? (8'h9f) : (8'hb5))) ? (((8'hb8) ? (8'ha0) : (8'hb2)) & ((8'ha2) - (7'h42))) : (((8'h9d) ? (8'haa) : (8'hbd)) - (|(7'h40))))) ? {(~^(|((8'hb2) ? (8'hba) : (8'hb7))))} : {(&(~|(-(8'ha9)))), (((^~(8'hab)) >= (8'hbd)) <<< (((8'ha9) ? (8'hab) : (8'hba)) <<< ((7'h40) ? (8'haa) : (8'ha8))))}))
(y, clk, wire54, wire53, wire52, wire51, wire50);
  output wire [(32'he9):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire54;
  input wire signed [(4'hb):(1'h0)] wire53;
  input wire signed [(5'h10):(1'h0)] wire52;
  input wire [(5'h14):(1'h0)] wire51;
  input wire [(5'h12):(1'h0)] wire50;
  wire [(3'h4):(1'h0)] wire75;
  wire signed [(5'h14):(1'h0)] wire74;
  wire signed [(5'h13):(1'h0)] wire73;
  wire signed [(2'h2):(1'h0)] wire69;
  wire signed [(3'h5):(1'h0)] wire68;
  wire [(3'h5):(1'h0)] wire67;
  wire [(3'h5):(1'h0)] wire63;
  wire signed [(4'hf):(1'h0)] wire62;
  wire signed [(5'h14):(1'h0)] wire61;
  wire signed [(4'hd):(1'h0)] wire60;
  wire signed [(4'h8):(1'h0)] wire59;
  wire signed [(4'hf):(1'h0)] wire58;
  wire signed [(5'h13):(1'h0)] wire57;
  wire [(4'h9):(1'h0)] wire56;
  wire [(2'h3):(1'h0)] wire55;
  reg [(4'ha):(1'h0)] reg72 = (1'h0);
  reg [(4'h8):(1'h0)] reg71 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg70 = (1'h0);
  reg [(4'ha):(1'h0)] reg66 = (1'h0);
  reg [(5'h11):(1'h0)] reg65 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg64 = (1'h0);
  assign y = {wire75,
                 wire74,
                 wire73,
                 wire69,
                 wire68,
                 wire67,
                 wire63,
                 wire62,
                 wire61,
                 wire60,
                 wire59,
                 wire58,
                 wire57,
                 wire56,
                 wire55,
                 reg72,
                 reg71,
                 reg70,
                 reg66,
                 reg65,
                 reg64,
                 (1'h0)};
  assign wire55 = wire51[(2'h2):(2'h2)];
  assign wire56 = $unsigned((~|($unsigned({wire50}) << wire55)));
  assign wire57 = wire55;
  assign wire58 = wire51[(3'h4):(1'h0)];
  assign wire59 = ($signed(wire56) == $signed((wire57[(4'hc):(4'h8)] ?
                      (8'ha9) : $signed($signed(wire50)))));
  assign wire60 = wire51[(5'h14):(5'h10)];
  assign wire61 = $unsigned((-wire58));
  assign wire62 = wire51[(4'hb):(2'h3)];
  assign wire63 = $unsigned((-wire59[(3'h5):(1'h0)]));
  always
    @(posedge clk) begin
      reg64 <= $signed($unsigned((({wire55} ?
          wire63 : wire60[(3'h4):(2'h2)]) == wire53[(3'h6):(1'h1)])));
      reg65 <= wire50[(3'h7):(3'h5)];
      reg66 <= {$unsigned($signed($signed(wire55[(1'h0):(1'h0)]))),
          ((-$signed((wire55 * wire54))) ?
              {(wire58[(3'h6):(2'h2)] ?
                      (wire50 ?
                          wire61 : wire51) : $unsigned(wire61))} : ((wire59 ?
                      wire58 : $unsigned(reg65)) ?
                  wire56 : (wire56[(3'h7):(3'h5)] ?
                      (wire60 ? wire50 : (8'hb0)) : (8'ha2))))};
    end
  assign wire67 = wire62;
  assign wire68 = (-wire55[(1'h0):(1'h0)]);
  assign wire69 = (8'hb8);
  always
    @(posedge clk) begin
      reg70 <= $signed({wire63[(2'h3):(2'h2)],
          ((8'haa) > ((&wire56) ? (reg66 <= reg65) : wire58))});
      reg71 <= $signed((~&((wire69[(2'h2):(1'h0)] ?
          wire50[(2'h2):(1'h0)] : (wire51 == wire52)) <= $unsigned($unsigned(wire58)))));
      reg72 <= ($signed(((reg70 == (wire53 + wire62)) ?
          ((wire69 ? wire62 : wire57) ?
              (~^wire50) : $unsigned(wire62)) : $signed((~^wire52)))) && $unsigned($unsigned($unsigned(wire51))));
    end
  assign wire73 = (|$signed((&(~|(wire54 ? wire56 : wire61)))));
  assign wire74 = (~&reg66[(3'h6):(3'h5)]);
  assign wire75 = $unsigned({reg64[(2'h2):(2'h2)]});
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module246
#(parameter param258 = (((&((!(8'ha3)) ? (8'h9f) : ((8'hbd) ? (8'hba) : (7'h44)))) * {(((8'hb3) << (8'ha7)) ? ((8'hb5) || (8'hb5)) : (8'hb5))}) ? (((((8'ha2) * (8'ha5)) + {(8'h9d)}) ? (((8'hb4) + (8'h9f)) ? ((8'ha4) & (8'ha1)) : ((8'h9c) ? (8'hb7) : (8'hbd))) : (((8'ha3) & (8'haf)) < {(7'h43), (8'hbe)})) ? (((7'h40) ? ((8'ha2) * (8'ha6)) : {(7'h43), (7'h44)}) ? (~^(^~(8'hb5))) : (|{(7'h41)})) : ((+(&(8'hb2))) ? (&(&(8'hb0))) : ((8'hb9) ? ((8'hae) ^~ (8'hb5)) : ((8'haa) ? (8'ha3) : (8'hb0))))) : ((((&(7'h40)) ? ((8'ha0) - (8'h9e)) : (~(7'h43))) <= {((7'h40) ? (8'hab) : (8'hb1))}) - ((((8'hbb) + (7'h40)) ? {(8'hbc)} : ((8'ha3) ? (7'h40) : (8'hbe))) ? {((7'h42) <<< (8'hae)), (~|(7'h42))} : {{(8'had), (8'h9c)}, (~(8'hb4))}))), 
parameter param259 = {(((^~(^~param258)) ? ((&param258) ? (8'hb2) : (param258 ? param258 : param258)) : (!(param258 ? param258 : param258))) & (((&param258) ? param258 : (|param258)) <= param258))})
(y, clk, wire251, wire250, wire249, wire248, wire247);
  output wire [(32'h47):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hf):(1'h0)] wire251;
  input wire signed [(5'h10):(1'h0)] wire250;
  input wire signed [(5'h11):(1'h0)] wire249;
  input wire [(4'hc):(1'h0)] wire248;
  input wire [(4'h9):(1'h0)] wire247;
  wire [(4'hb):(1'h0)] wire257;
  wire signed [(3'h4):(1'h0)] wire256;
  wire signed [(5'h14):(1'h0)] wire255;
  wire [(4'hb):(1'h0)] wire254;
  wire [(4'hd):(1'h0)] wire253;
  wire [(4'hb):(1'h0)] wire252;
  assign y = {wire257, wire256, wire255, wire254, wire253, wire252, (1'h0)};
  assign wire252 = {(wire248 ?
                           wire251[(3'h5):(2'h2)] : ($signed(wire249) >= wire248)),
                       $signed(wire250[(4'hb):(1'h0)])};
  assign wire253 = $signed($signed((wire251 && $signed(wire249))));
  assign wire254 = {$signed((+$unsigned(wire251))), wire250};
  assign wire255 = {wire249[(4'hf):(3'h4)]};
  assign wire256 = (8'h9f);
  assign wire257 = (^~wire251);
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module186
#(parameter param241 = (({((^(8'hae)) == {(8'hb1)}), (8'h9e)} ? ((^~(^~(8'hb8))) <<< (((8'hb9) ? (8'hb7) : (8'haa)) ~^ ((8'hb9) & (7'h42)))) : (&{(~^(8'ha1))})) > {(7'h42), (&((8'hb0) <<< ((8'h9c) ? (7'h43) : (7'h40))))}))
(y, clk, wire190, wire189, wire188, wire187);
  output wire [(32'h226):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h6):(1'h0)] wire190;
  input wire signed [(3'h6):(1'h0)] wire189;
  input wire [(5'h12):(1'h0)] wire188;
  input wire signed [(5'h12):(1'h0)] wire187;
  wire [(4'hd):(1'h0)] wire240;
  wire signed [(5'h13):(1'h0)] wire239;
  wire signed [(3'h6):(1'h0)] wire238;
  wire signed [(3'h6):(1'h0)] wire236;
  wire signed [(4'hd):(1'h0)] wire235;
  wire signed [(3'h4):(1'h0)] wire234;
  wire [(4'hc):(1'h0)] wire233;
  wire signed [(3'h6):(1'h0)] wire232;
  wire [(5'h10):(1'h0)] wire223;
  wire [(4'hc):(1'h0)] wire222;
  wire [(3'h4):(1'h0)] wire215;
  wire signed [(5'h12):(1'h0)] wire214;
  wire signed [(3'h7):(1'h0)] wire213;
  wire [(4'hb):(1'h0)] wire196;
  wire signed [(2'h3):(1'h0)] wire195;
  wire [(4'hb):(1'h0)] wire194;
  wire signed [(5'h10):(1'h0)] wire191;
  reg signed [(3'h5):(1'h0)] reg237 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg231 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg230 = (1'h0);
  reg [(4'ha):(1'h0)] reg227 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg226 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg225 = (1'h0);
  reg [(4'h9):(1'h0)] reg224 = (1'h0);
  reg [(4'ha):(1'h0)] reg221 = (1'h0);
  reg [(3'h4):(1'h0)] reg219 = (1'h0);
  reg [(5'h10):(1'h0)] reg218 = (1'h0);
  reg [(2'h2):(1'h0)] reg217 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg216 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg211 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg208 = (1'h0);
  reg [(5'h14):(1'h0)] reg207 = (1'h0);
  reg [(5'h13):(1'h0)] reg204 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg203 = (1'h0);
  reg [(4'hb):(1'h0)] reg202 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg200 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg199 = (1'h0);
  reg [(5'h15):(1'h0)] reg193 = (1'h0);
  reg [(4'hc):(1'h0)] reg192 = (1'h0);
  reg [(4'h8):(1'h0)] forvar229 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg228 = (1'h0);
  reg [(5'h11):(1'h0)] forvar220 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg212 = (1'h0);
  reg [(5'h10):(1'h0)] reg210 = (1'h0);
  reg [(4'hf):(1'h0)] forvar209 = (1'h0);
  reg [(4'h8):(1'h0)] reg206 = (1'h0);
  reg [(3'h7):(1'h0)] forvar205 = (1'h0);
  reg [(2'h2):(1'h0)] reg201 = (1'h0);
  reg [(5'h10):(1'h0)] forvar198 = (1'h0);
  reg [(2'h2):(1'h0)] forvar197 = (1'h0);
  assign y = {wire240,
                 wire239,
                 wire238,
                 wire236,
                 wire235,
                 wire234,
                 wire233,
                 wire232,
                 wire223,
                 wire222,
                 wire215,
                 wire214,
                 wire213,
                 wire196,
                 wire195,
                 wire194,
                 wire191,
                 reg237,
                 reg231,
                 reg230,
                 reg227,
                 reg226,
                 reg225,
                 reg224,
                 reg221,
                 reg219,
                 reg218,
                 reg217,
                 reg216,
                 reg211,
                 reg208,
                 reg207,
                 reg204,
                 reg203,
                 reg202,
                 reg200,
                 reg199,
                 reg193,
                 reg192,
                 forvar229,
                 reg228,
                 forvar220,
                 reg212,
                 reg210,
                 forvar209,
                 reg206,
                 forvar205,
                 reg201,
                 forvar198,
                 forvar197,
                 (1'h0)};
  assign wire191 = $signed({(((8'hbb) < $signed(wire189)) >>> $unsigned($signed(wire189))),
                       (~^(+(wire189 ? wire190 : (7'h41))))});
  always
    @(posedge clk) begin
      reg192 <= wire188[(3'h6):(1'h0)];
      reg193 <= wire188;
    end
  assign wire194 = $signed(($unsigned(wire187) ?
                       (-wire189[(2'h2):(2'h2)]) : ($unsigned((wire190 - (8'hba))) ?
                           $unsigned((wire191 ?
                               wire189 : wire190)) : ((~|wire191) ?
                               reg193 : wire189[(2'h3):(1'h1)]))));
  assign wire195 = $unsigned($unsigned(($signed(((8'hb1) ? (8'haf) : wire190)) ?
                       ((-wire188) - $unsigned(wire191)) : wire190)));
  assign wire196 = ((+$unsigned(reg193)) <= {((~^(^reg193)) >= (~|(wire190 || wire188)))});
  always
    @(posedge clk) begin
      for (forvar197 = (1'h0); (forvar197 < (3'h4)); forvar197 = (forvar197 + (1'h1)))
        begin
          for (forvar198 = (1'h0); (forvar198 < (3'h4)); forvar198 = (forvar198 + (1'h1)))
            begin
              reg199 <= wire195;
              reg200 <= forvar197[(1'h0):(1'h0)];
              reg201 = (wire187[(3'h5):(3'h4)] ?
                  reg193[(5'h14):(4'hb)] : (~|reg199[(2'h3):(1'h1)]));
              reg202 <= $signed((((((8'h9d) ? wire190 : wire187) ?
                      reg201[(1'h0):(1'h0)] : (wire191 + wire190)) - (&$unsigned((8'hbc)))) ?
                  $unsigned($signed((wire189 ?
                      (7'h43) : wire188))) : $signed($unsigned($unsigned((8'had))))));
              reg203 <= wire190;
            end
          reg204 <= {(~^(^(wire190 ? wire188[(3'h7):(3'h5)] : forvar197)))};
        end
      for (forvar205 = (1'h0); (forvar205 < (1'h0)); forvar205 = (forvar205 + (1'h1)))
        begin
          reg206 = {forvar198, (~(+{(wire195 >>> reg201)}))};
          reg207 <= (&($unsigned($signed((forvar205 > wire190))) ?
              ($signed({wire190,
                  forvar205}) && ((~^reg199) * wire196)) : wire187));
        end
      reg208 <= reg199;
      for (forvar209 = (1'h0); (forvar209 < (1'h0)); forvar209 = (forvar209 + (1'h1)))
        begin
          reg210 = (|reg204);
          reg211 <= (wire187 ? reg208 : wire191);
          reg212 = (forvar205[(2'h2):(2'h2)] ? (7'h40) : reg192);
        end
    end
  assign wire213 = (~$unsigned($unsigned({(wire196 ? reg202 : reg202)})));
  assign wire214 = ({$unsigned((~(|(8'hb0))))} < $signed({(!(~^reg208)),
                       ($signed((8'hb5)) > $signed(reg211))}));
  assign wire215 = (^wire191[(4'h9):(2'h3)]);
  always
    @(posedge clk) begin
      reg216 <= $signed((~|{$unsigned((wire215 ? reg204 : reg192)),
          ((^wire194) ?
              ((8'ha7) ? wire191 : (7'h40)) : reg208[(4'hb):(4'h8)])}));
      reg217 <= wire189;
      reg218 <= (wire195 ^ $signed({({reg203} ?
              (wire195 ~^ wire190) : reg199[(3'h5):(2'h2)])}));
      reg219 <= reg218;
      for (forvar220 = (1'h0); (forvar220 < (1'h1)); forvar220 = (forvar220 + (1'h1)))
        begin
          reg221 <= $unsigned($unsigned((forvar220 == $signed($signed(reg203)))));
        end
    end
  assign wire222 = (reg202 + {(((~&reg200) ?
                               reg221[(4'h8):(3'h5)] : wire190[(1'h0):(1'h0)]) ?
                           reg193[(2'h3):(1'h1)] : reg208),
                       (8'h9e)});
  assign wire223 = (~&{{reg192[(3'h7):(3'h6)]}});
  always
    @(posedge clk) begin
      reg224 <= (reg217 + {($unsigned(wire187) > (^(8'haa))), reg218});
      reg225 <= $signed(reg208);
    end
  always
    @(posedge clk) begin
      reg226 <= (wire222 ?
          wire194[(2'h3):(2'h3)] : (((reg204[(4'he):(4'ha)] | {wire223}) ~^ ((wire196 > reg204) ?
              (wire189 | reg221) : (wire194 ?
                  wire222 : (8'ha3)))) >> (|(8'hac))));
      reg227 <= (|((({reg202} >>> $unsigned(reg203)) ?
              (wire223[(4'hb):(3'h4)] ?
                  (~|reg192) : $signed(reg221)) : wire191[(1'h1):(1'h1)]) ?
          (~|$unsigned(reg218)) : $signed(reg199)));
      reg228 = wire214[(4'hb):(3'h7)];
      for (forvar229 = (1'h0); (forvar229 < (1'h1)); forvar229 = (forvar229 + (1'h1)))
        begin
          reg230 <= (((&((-reg227) ? (-reg202) : $signed(forvar229))) ?
              ($unsigned((wire195 ?
                  wire191 : reg227)) - wire190) : (!((~|wire194) < (+reg216)))) >= (~(reg200 ?
              $signed($unsigned(reg218)) : (((8'hb4) ?
                  reg217 : reg224) ~^ (reg219 & reg204)))));
        end
      reg231 <= $unsigned($signed({(|$signed(reg217)), (!(wire194 | reg192))}));
    end
  assign wire232 = {$unsigned((reg219[(1'h0):(1'h0)] + ($unsigned(reg231) ?
                           (reg218 ? (8'h9d) : reg199) : (reg203 || wire188)))),
                       reg224[(3'h5):(3'h4)]};
  assign wire233 = reg224[(3'h4):(2'h3)];
  assign wire234 = $signed($unsigned(((^~reg226) ?
                       reg227[(4'h8):(4'h8)] : ((&wire194) & (reg208 ^ reg202)))));
  assign wire235 = reg225;
  assign wire236 = ((^~wire233) ?
                       $signed((~reg217[(2'h2):(2'h2)])) : $unsigned($signed((+{wire194,
                           reg192}))));
  always
    @(posedge clk) begin
      reg237 <= $signed(reg199);
    end
  assign wire238 = (8'hab);
  assign wire239 = reg200;
  assign wire240 = (wire190 ?
                       reg199[(3'h6):(3'h4)] : $unsigned(($unsigned((^(8'hbc))) ?
                           reg199 : $unsigned({wire191}))));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module173
#(parameter param183 = ((~&((^((8'ha7) > (8'hb9))) ^~ (((8'h9f) ? (8'h9c) : (7'h40)) ? {(8'ha8), (8'ha0)} : {(8'hbb), (8'haa)}))) || (+{(((8'ha5) ? (8'ha8) : (8'hb2)) >>> ((8'hb0) <= (7'h40))), (7'h42)})))
(y, clk, wire178, wire177, wire176, wire175, wire174);
  output wire [(32'h22):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire178;
  input wire signed [(5'h14):(1'h0)] wire177;
  input wire [(4'h9):(1'h0)] wire176;
  input wire signed [(3'h7):(1'h0)] wire175;
  input wire signed [(4'hf):(1'h0)] wire174;
  wire [(4'ha):(1'h0)] wire182;
  wire signed [(2'h3):(1'h0)] wire181;
  wire signed [(4'h8):(1'h0)] wire180;
  wire [(4'hc):(1'h0)] wire179;
  assign y = {wire182, wire181, wire180, wire179, (1'h0)};
  assign wire179 = ({(((wire174 ^ wire178) ? (&wire178) : (~|(8'hbc))) ?
                               $signed((wire177 ?
                                   wire174 : wire175)) : $unsigned((wire177 | wire175))),
                           ($unsigned((wire175 < wire175)) ?
                               wire177[(4'h8):(3'h4)] : wire178)} ?
                       wire177 : ((8'hb7) ?
                           $signed($unsigned((8'hb9))) : ($unsigned(((8'ha8) ?
                                   (8'h9d) : wire177)) ?
                               $unsigned($signed((8'hbb))) : ((wire177 > wire178) != (wire174 ?
                                   wire176 : wire174)))));
  assign wire180 = $signed((~((~(-wire175)) ?
                       $signed((^~wire175)) : $signed(wire177[(4'hd):(4'h8)]))));
  assign wire181 = wire180;
  assign wire182 = $unsigned((~&$unsigned($signed((|wire175)))));
endmodule