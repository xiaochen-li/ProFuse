(* use_dsp48="no" *) (* use_dsp="no" *) module top  (y, clk, wire0, wire1, wire2, wire3);
  output wire [(32'h59d):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(3'h7):(1'h0)] wire0;
  input wire [(4'hd):(1'h0)] wire1;
  input wire [(2'h2):(1'h0)] wire2;
  input wire [(5'h15):(1'h0)] wire3;
  wire [(4'h9):(1'h0)] wire691;
  wire signed [(5'h10):(1'h0)] wire690;
  wire [(4'hc):(1'h0)] wire4;
  wire [(2'h3):(1'h0)] wire70;
  wire [(5'h12):(1'h0)] wire71;
  wire signed [(3'h7):(1'h0)] wire461;
  wire signed [(3'h6):(1'h0)] wire670;
  reg [(5'h11):(1'h0)] reg719 = (1'h0);
  reg [(5'h11):(1'h0)] reg718 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg713 = (1'h0);
  reg [(4'h9):(1'h0)] reg711 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg709 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg708 = (1'h0);
  reg [(3'h6):(1'h0)] reg707 = (1'h0);
  reg [(5'h12):(1'h0)] reg704 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg702 = (1'h0);
  reg [(3'h6):(1'h0)] reg701 = (1'h0);
  reg [(3'h7):(1'h0)] reg699 = (1'h0);
  reg [(2'h3):(1'h0)] reg698 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg697 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg694 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg693 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg689 = (1'h0);
  reg [(4'hc):(1'h0)] reg687 = (1'h0);
  reg [(4'h9):(1'h0)] reg683 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg676 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg674 = (1'h0);
  reg [(4'hd):(1'h0)] reg672 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg6 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg8 = (1'h0);
  reg [(2'h2):(1'h0)] reg10 = (1'h0);
  reg [(4'h8):(1'h0)] reg11 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg12 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg15 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg17 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg18 = (1'h0);
  reg [(4'hd):(1'h0)] reg22 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg23 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg24 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg26 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg19 = (1'h0);
  reg [(4'he):(1'h0)] reg29 = (1'h0);
  reg [(4'hc):(1'h0)] reg30 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg31 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg34 = (1'h0);
  reg [(4'he):(1'h0)] reg36 = (1'h0);
  reg [(5'h11):(1'h0)] reg38 = (1'h0);
  reg [(4'hd):(1'h0)] reg39 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg41 = (1'h0);
  reg [(5'h14):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg43 = (1'h0);
  reg [(3'h5):(1'h0)] reg49 = (1'h0);
  reg [(3'h6):(1'h0)] reg51 = (1'h0);
  reg [(4'h9):(1'h0)] reg52 = (1'h0);
  reg [(4'he):(1'h0)] reg54 = (1'h0);
  reg [(5'h10):(1'h0)] reg55 = (1'h0);
  reg [(4'hd):(1'h0)] reg56 = (1'h0);
  reg signed [(4'he):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg58 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg59 = (1'h0);
  reg [(4'ha):(1'h0)] reg61 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg63 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg65 = (1'h0);
  reg [(5'h10):(1'h0)] reg66 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg69 = (1'h0);
  reg [(4'hd):(1'h0)] reg717 = (1'h0);
  reg [(4'hd):(1'h0)] reg716 = (1'h0);
  reg [(5'h15):(1'h0)] reg715 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar714 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg712 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar710 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg706 = (1'h0);
  reg [(5'h11):(1'h0)] reg705 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg703 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg700 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar696 = (1'h0);
  reg [(5'h12):(1'h0)] reg695 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar692 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg688 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg686 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg685 = (1'h0);
  reg [(5'h13):(1'h0)] reg684 = (1'h0);
  reg [(4'hd):(1'h0)] reg682 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg681 = (1'h0);
  reg [(4'hc):(1'h0)] reg680 = (1'h0);
  reg [(3'h6):(1'h0)] reg679 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg678 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg673 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg677 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg675 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar673 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg68 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg67 = (1'h0);
  reg [(5'h12):(1'h0)] forvar64 = (1'h0);
  reg [(4'hb):(1'h0)] reg62 = (1'h0);
  reg [(5'h14):(1'h0)] reg60 = (1'h0);
  reg [(3'h7):(1'h0)] reg53 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar53 = (1'h0);
  reg [(4'hc):(1'h0)] reg50 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar48 = (1'h0);
  reg signed [(4'he):(1'h0)] reg47 = (1'h0);
  reg [(4'he):(1'h0)] reg46 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar45 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg44 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar40 = (1'h0);
  reg [(5'h15):(1'h0)] reg37 = (1'h0);
  reg [(4'he):(1'h0)] reg35 = (1'h0);
  reg [(3'h6):(1'h0)] reg33 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg32 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg28 = (1'h0);
  reg [(3'h7):(1'h0)] forvar27 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar23 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg25 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg21 = (1'h0);
  reg [(5'h13):(1'h0)] reg20 = (1'h0);
  reg [(4'hd):(1'h0)] forvar19 = (1'h0);
  reg [(2'h3):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar14 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg13 = (1'h0);
  reg [(3'h4):(1'h0)] forvar10 = (1'h0);
  reg [(4'hd):(1'h0)] reg9 = (1'h0);
  reg [(4'hc):(1'h0)] forvar7 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg5 = (1'h0);
  assign y = {wire691,
                 wire690,
                 wire4,
                 wire70,
                 wire71,
                 wire461,
                 wire670,
                 reg719,
                 reg718,
                 reg713,
                 reg711,
                 reg709,
                 reg708,
                 reg707,
                 reg704,
                 reg702,
                 reg701,
                 reg699,
                 reg698,
                 reg697,
                 reg694,
                 reg693,
                 reg689,
                 reg687,
                 reg683,
                 reg676,
                 reg674,
                 reg672,
                 reg6,
                 reg8,
                 reg10,
                 reg11,
                 reg12,
                 reg15,
                 reg17,
                 reg18,
                 reg22,
                 reg23,
                 reg24,
                 reg26,
                 reg19,
                 reg29,
                 reg30,
                 reg31,
                 reg34,
                 reg36,
                 reg38,
                 reg39,
                 reg41,
                 reg42,
                 reg43,
                 reg49,
                 reg51,
                 reg52,
                 reg54,
                 reg55,
                 reg56,
                 reg57,
                 reg58,
                 reg59,
                 reg61,
                 reg63,
                 reg65,
                 reg66,
                 reg69,
                 reg717,
                 reg716,
                 reg715,
                 forvar714,
                 reg712,
                 forvar710,
                 reg706,
                 reg705,
                 reg703,
                 reg700,
                 forvar696,
                 reg695,
                 forvar692,
                 reg688,
                 reg686,
                 reg685,
                 reg684,
                 reg682,
                 reg681,
                 reg680,
                 reg679,
                 reg678,
                 reg673,
                 reg677,
                 reg675,
                 forvar673,
                 reg68,
                 reg67,
                 forvar64,
                 reg62,
                 reg60,
                 reg53,
                 forvar53,
                 reg50,
                 forvar48,
                 reg47,
                 reg46,
                 forvar45,
                 reg44,
                 forvar40,
                 reg37,
                 reg35,
                 reg33,
                 reg32,
                 reg28,
                 forvar27,
                 forvar23,
                 reg25,
                 reg21,
                 reg20,
                 forvar19,
                 reg16,
                 forvar14,
                 reg13,
                 forvar10,
                 reg9,
                 forvar7,
                 reg5,
                 (1'h0)};
  assign wire4 = $signed(wire3[(5'h14):(4'hf)]);
  always
    @(posedge clk) begin
      if ($signed((8'ha3)))
        begin
          reg5 = ((($signed((wire3 < wire4)) || $unsigned($unsigned(wire1))) ?
              ((!(wire4 >> wire4)) ?
                  wire0 : (!((7'h43) >> wire1))) : wire1) > $unsigned((wire3 ?
              (~|wire2[(1'h1):(1'h1)]) : $unsigned($unsigned(wire4)))));
        end
      else
        begin
          reg5 = ((+(^~$unsigned(wire2))) ? reg5[(3'h7):(3'h4)] : wire4);
          reg6 <= (&$unsigned(($unsigned(((8'hb1) ?
              wire3 : wire0)) > (((8'hbb) ? wire0 : wire0) ?
              (~^wire0) : ((8'hb3) <= wire0)))));
          for (forvar7 = (1'h0); (forvar7 < (3'h4)); forvar7 = (forvar7 + (1'h1)))
            begin
              reg8 <= {$unsigned((wire4 || ($signed(wire0) ?
                      $signed(wire3) : ((8'hbf) >= reg5))))};
              reg9 = ((7'h41) ^ wire2[(1'h0):(1'h0)]);
            end
        end
    end
  always
    @(posedge clk) begin
      if ((wire1[(3'h5):(2'h3)] << ((8'hb7) ?
          wire2[(2'h2):(1'h0)] : ((~(wire1 == wire4)) ?
              {$unsigned(wire4)} : $signed((reg6 ? wire0 : wire4))))))
        begin
          reg10 <= (reg6[(1'h1):(1'h0)] ~^ {{wire1},
              $unsigned(wire3[(5'h10):(4'hd)])});
          reg11 <= (~|($signed((&reg10[(1'h1):(1'h0)])) > (&reg8)));
        end
      else
        begin
          for (forvar10 = (1'h0); (forvar10 < (2'h2)); forvar10 = (forvar10 + (1'h1)))
            begin
              reg11 <= (((&(7'h40)) < (wire3[(5'h15):(3'h7)] ~^ $unsigned($signed(reg10)))) ?
                  reg6 : $signed((reg8 | wire2)));
            end
          reg12 <= $unsigned(reg6);
          reg13 = (^{reg10, (reg8 == reg8[(4'he):(2'h3)])});
          for (forvar14 = (1'h0); (forvar14 < (1'h0)); forvar14 = (forvar14 + (1'h1)))
            begin
              reg15 <= (reg6[(3'h7):(3'h7)] ?
                  $unsigned(((|(reg8 ? wire2 : (8'hbf))) ?
                      $unsigned($unsigned(wire1)) : $unsigned((wire4 ?
                          wire0 : (8'hb3))))) : (|reg8));
              reg16 = ($unsigned((forvar10[(1'h0):(1'h0)] != wire1[(3'h4):(2'h2)])) + $signed($unsigned(($signed((8'ha0)) ?
                  reg12 : $signed(reg15)))));
            end
        end
      reg17 <= (-{($unsigned((+wire2)) ?
              (^~(reg16 ? reg8 : (7'h43))) : {$unsigned(reg15)})});
    end
  always
    @(posedge clk) begin
      if (wire4)
        begin
          reg18 <= $signed($signed(wire1[(3'h7):(3'h5)]));
          for (forvar19 = (1'h0); (forvar19 < (3'h4)); forvar19 = (forvar19 + (1'h1)))
            begin
              reg20 = (((-(~&wire0)) ^ reg15[(3'h4):(1'h0)]) ?
                  (reg11 ^ (^~(8'hb4))) : $unsigned($unsigned((+forvar19))));
              reg21 = (8'hba);
            end
          if ((($signed($unsigned({wire1})) >> $unsigned($unsigned(reg6[(4'hb):(1'h0)]))) << $signed((reg11 + (&reg21)))))
            begin
              reg22 <= (8'hbb);
              reg23 <= ((^~((reg22 ^ wire2) >= ((wire4 < reg12) ?
                  (~^forvar19) : $unsigned(reg22)))) >> ({((8'h9e) ~^ (wire4 ?
                          wire0 : reg8))} ?
                  {((reg22 - reg6) ?
                          $unsigned(wire3) : $unsigned(reg11))} : (($signed(reg6) ?
                          reg11 : $unsigned(reg15)) ?
                      reg8 : (8'hb4))));
              reg24 <= ($unsigned((~&reg12)) ?
                  (8'hb8) : (reg6[(4'hc):(4'hb)] ?
                      wire3[(3'h7):(2'h2)] : {{$unsigned(reg17), (8'hb4)},
                          $unsigned((~|reg15))}));
            end
          else
            begin
              reg22 <= $unsigned($signed(((reg17[(3'h6):(1'h0)] ?
                  $unsigned((8'h9f)) : reg10[(1'h1):(1'h1)]) >= ((wire3 <= reg8) ?
                  (+wire3) : reg10[(1'h1):(1'h1)]))));
              reg23 <= (((wire0 <<< $unsigned(wire1)) + reg18) ?
                  $unsigned($unsigned((^~$unsigned((8'hb4))))) : reg23[(4'hf):(3'h4)]);
              reg25 = {reg20};
              reg26 <= reg10;
            end
        end
      else
        begin
          reg18 <= {$unsigned(reg10),
              ({$signed(reg12)} ?
                  (^~(+(wire2 ?
                      forvar19 : reg24))) : $signed(wire3[(1'h1):(1'h1)]))};
          reg19 <= reg21;
          reg22 <= reg20[(1'h1):(1'h1)];
          for (forvar23 = (1'h0); (forvar23 < (1'h0)); forvar23 = (forvar23 + (1'h1)))
            begin
              reg24 <= ((reg26 << forvar23[(2'h2):(1'h0)]) ?
                  $unsigned((&$signed($signed(wire4)))) : ($signed(reg15) < $unsigned(((reg10 ?
                          (8'hb2) : (8'haa)) ?
                      (reg19 >> reg8) : reg22))));
              reg26 <= $unsigned((+(~wire4)));
            end
        end
      for (forvar27 = (1'h0); (forvar27 < (1'h1)); forvar27 = (forvar27 + (1'h1)))
        begin
          reg28 = ((7'h41) ? $unsigned($unsigned(forvar23)) : reg15);
        end
      reg29 <= (~^(reg11[(3'h5):(1'h1)] ?
          (($unsigned(reg19) >>> reg19[(4'hf):(4'he)]) ?
              (wire2 ? wire2 : $unsigned(reg15)) : ((wire4 <= reg19) ?
                  ((7'h43) >= reg10) : $unsigned(wire2))) : (~^$signed($signed(reg17)))));
      reg30 <= (8'hb4);
    end
  always
    @(posedge clk) begin
      reg31 <= reg15;
      reg32 = wire2[(1'h1):(1'h0)];
      reg33 = $unsigned($unsigned(reg29));
    end
  always
    @(posedge clk) begin
      reg34 <= wire2[(1'h0):(1'h0)];
      reg35 = {((({reg26, wire3} & {reg11, reg12}) | reg29) ?
              $unsigned(((reg17 ? reg31 : reg23) ?
                  (-reg22) : (reg10 ?
                      reg17 : reg22))) : ($signed($signed((8'ha3))) ?
                  ((|reg6) ?
                      $unsigned(wire1) : $signed(wire3)) : $unsigned((reg11 < (8'haa))))),
          $signed(reg12[(2'h2):(1'h0)])};
      reg36 <= ((~|reg10[(2'h2):(2'h2)]) & (reg31[(1'h0):(1'h0)] ?
          reg31 : wire3));
    end
  always
    @(posedge clk) begin
      reg37 = ((reg10[(1'h1):(1'h0)] ?
          ($unsigned($signed(reg34)) ?
              ((8'hbd) & $signed(reg29)) : ({reg10,
                  reg11} < (7'h42))) : wire1[(3'h7):(1'h1)]) & reg6[(4'hb):(3'h7)]);
      reg38 <= $signed(reg6);
      reg39 <= $unsigned(reg23);
      for (forvar40 = (1'h0); (forvar40 < (1'h1)); forvar40 = (forvar40 + (1'h1)))
        begin
          reg41 <= $unsigned($unsigned($signed({$unsigned((8'hbe))})));
          reg42 <= reg26;
          reg43 <= {(7'h43),
              $signed($unsigned(((reg26 * (8'hbe)) ?
                  wire0[(3'h6):(1'h0)] : $unsigned(reg30))))};
        end
    end
  always
    @(posedge clk) begin
      reg44 = wire4[(3'h6):(2'h2)];
      for (forvar45 = (1'h0); (forvar45 < (2'h3)); forvar45 = (forvar45 + (1'h1)))
        begin
          reg46 = ((^~(+$signed((reg22 ? reg42 : (8'h9d))))) ?
              ($signed((~^(reg38 ? (8'hb0) : (8'hbe)))) ?
                  $unsigned(reg15) : $unsigned((wire1 ?
                      {reg34, (8'hbe)} : {reg26,
                          wire3}))) : ((^~reg38[(4'ha):(2'h2)]) ?
                  ((^~(reg31 ~^ forvar45)) ?
                      reg10 : wire4) : wire2[(1'h0):(1'h0)]));
          reg47 = {$unsigned(reg11[(3'h4):(2'h2)]), (~reg6)};
          for (forvar48 = (1'h0); (forvar48 < (3'h4)); forvar48 = (forvar48 + (1'h1)))
            begin
              reg49 <= reg44;
              reg50 = reg18;
              reg51 <= $signed(reg15);
              reg52 <= ($signed(($unsigned((8'hbb)) >= $signed((reg29 ?
                  reg39 : (8'hb8))))) ^ ((reg51[(1'h0):(1'h0)] ^ (~|(reg34 << reg31))) - (8'hb3)));
            end
        end
      if (reg29[(4'ha):(3'h7)])
        begin
          for (forvar53 = (1'h0); (forvar53 < (2'h3)); forvar53 = (forvar53 + (1'h1)))
            begin
              reg54 <= {(reg22[(2'h2):(1'h0)] ?
                      (~|reg49) : ($unsigned((wire0 * reg39)) ?
                          $unsigned((wire0 * reg17)) : reg46))};
              reg55 <= reg38;
              reg56 <= $signed(reg41[(4'h9):(3'h5)]);
              reg57 <= ((~&{wire3}) ?
                  (^(((forvar45 > reg42) == (reg43 ? reg39 : reg46)) ?
                      ((reg42 * reg43) ?
                          (|(8'ha3)) : (~|(8'hb7))) : $unsigned((^~reg47)))) : (|(forvar53[(4'h8):(3'h7)] > (+forvar53))));
            end
          reg58 <= reg49[(3'h4):(1'h1)];
        end
      else
        begin
          if ((~(8'hb0)))
            begin
              reg53 = wire0;
              reg54 <= $unsigned({({wire0} | ((reg24 ?
                      reg24 : reg49) >>> {reg52}))});
              reg55 <= wire4[(3'h5):(1'h0)];
              reg56 <= ((!reg43) ?
                  (reg31[(1'h1):(1'h1)] >= ($signed((reg43 != reg23)) | {(8'h9c),
                      (^reg52)})) : (({$unsigned(reg30)} > ((reg23 ?
                          reg43 : reg36) ?
                      {(8'hbe)} : $unsigned(reg53))) - (wire0 + reg22[(4'hd):(4'h8)])));
              reg57 <= ($signed((8'hba)) ?
                  (~|$signed($signed((reg8 ? wire4 : wire3)))) : (8'hbc));
            end
          else
            begin
              reg54 <= ((~^{$unsigned($signed(reg8)),
                      $signed((reg6 ? forvar53 : (7'h43)))}) ?
                  ($signed(reg18[(2'h3):(1'h0)]) ?
                      ((-reg42[(3'h5):(3'h5)]) ?
                          {(+reg43)} : ((|(8'ha1)) & (wire1 >> reg58))) : reg58) : (wire1[(4'h8):(2'h3)] != (~|((+(8'h9f)) < $unsigned(reg44)))));
              reg55 <= {reg57};
              reg56 <= reg11[(3'h7):(1'h1)];
              reg57 <= $signed(wire4[(3'h5):(3'h4)]);
              reg58 <= $signed($unsigned({reg31[(1'h1):(1'h1)],
                  ((^~reg18) + (|wire0))}));
            end
          if ((($unsigned((reg43 >> reg34[(5'h13):(3'h5)])) ^ $unsigned(((-reg47) ?
              reg29 : $unsigned(reg10)))) >>> ((reg46[(3'h4):(2'h3)] ?
              ((reg10 ? reg50 : (8'hb8)) ?
                  (reg19 >> wire1) : $signed(reg42)) : reg34) * $signed(wire2[(1'h1):(1'h1)]))))
            begin
              reg59 <= ($signed((reg57 ?
                      ((reg53 ?
                          wire0 : reg36) == reg54[(4'h9):(4'h9)]) : {{reg42},
                          (~|reg44)})) ?
                  $unsigned($signed($unsigned($unsigned(reg39)))) : reg46[(3'h6):(3'h5)]);
              reg60 = reg6[(4'hd):(2'h2)];
            end
          else
            begin
              reg59 <= wire2[(2'h2):(1'h0)];
              reg61 <= reg6[(4'hb):(4'ha)];
              reg62 = $unsigned($signed(reg50));
            end
          reg63 <= (~|($unsigned($unsigned($signed(reg10))) ?
              ((~&(-(8'hb3))) ?
                  reg29 : ($signed(wire4) <<< reg11[(3'h4):(2'h2)])) : reg49));
          for (forvar64 = (1'h0); (forvar64 < (1'h0)); forvar64 = (forvar64 + (1'h1)))
            begin
              reg65 <= (8'h9f);
              reg66 <= (~&$unsigned((+({reg11, forvar64} ?
                  reg46 : $unsigned(reg18)))));
              reg67 = ((~^reg24[(2'h2):(1'h1)]) ?
                  (((~&reg56[(4'hc):(4'h8)]) ~^ (~(reg55 ?
                      reg8 : reg6))) >> {$unsigned((~reg50)),
                      (reg56 ^~ reg46[(3'h6):(2'h3)])}) : {{reg47[(4'hb):(4'h8)]}});
              reg68 = $signed($signed($unsigned(((&reg65) ?
                  reg8[(1'h1):(1'h0)] : reg52))));
            end
        end
      reg69 <= $unsigned($signed(reg55[(4'hf):(4'hf)]));
    end
  assign wire70 = $signed(wire3);
  assign wire71 = (($unsigned(reg22) ? (8'hbc) : (8'hb2)) ^ ((8'hbe) ?
                      $signed((+(-reg65))) : (((8'ha5) ? reg61 : (8'hbc)) ?
                          (reg42 && $signed(reg55)) : (^~(~^wire2)))));
  module72 #() modinst462 (wire461, clk, reg12, reg43, reg6, reg57);
  module463 #() modinst671 (.clk(clk), .y(wire670), .wire467(wire1), .wire464(reg54), .wire465(reg22), .wire466(reg18));
  always
    @(posedge clk) begin
      reg672 <= wire3;
      if (reg31[(2'h2):(1'h1)])
        begin
          for (forvar673 = (1'h0); (forvar673 < (1'h1)); forvar673 = (forvar673 + (1'h1)))
            begin
              reg674 <= (+reg39[(3'h7):(3'h6)]);
              reg675 = (-(+(8'hb9)));
            end
          reg676 <= reg51[(1'h1):(1'h1)];
          reg677 = (reg8[(2'h3):(1'h0)] ~^ $unsigned(reg43[(3'h5):(1'h0)]));
        end
      else
        begin
          reg673 = reg29;
          if ($signed(reg30))
            begin
              reg675 = reg24;
              reg676 <= {$unsigned(reg63), (8'h9d)};
              reg677 = $unsigned(wire4);
              reg678 = reg42[(4'hc):(2'h3)];
              reg679 = ($signed((wire70[(1'h0):(1'h0)] << $signed((&(8'hbe))))) ?
                  $unsigned((reg52[(3'h5):(2'h2)] + ({reg49, (8'hb1)} ?
                      (reg66 ?
                          reg36 : (8'hbf)) : (wire4 == reg677)))) : ($signed(reg24) ^ $signed({wire670,
                      (^~reg56)})));
            end
          else
            begin
              reg674 <= $unsigned({$signed($signed(wire0))});
              reg675 = $unsigned(((((wire71 ? (8'ha2) : wire2) <<< (reg54 ?
                          reg52 : reg18)) ?
                      ($unsigned(reg49) ?
                          $signed(reg24) : (~&reg10)) : (-(8'ha5))) ?
                  (^($signed(reg42) ?
                      (&reg679) : $signed((8'hb8)))) : {{reg674},
                      (~(reg673 < wire670))}));
              reg677 = ($unsigned((reg42 && (reg24[(1'h1):(1'h1)] ?
                  reg675[(1'h0):(1'h0)] : $unsigned(reg677)))) * reg66[(3'h5):(3'h5)]);
            end
          reg680 = (reg26[(3'h6):(3'h6)] || $signed(({reg69} > (&$signed(reg52)))));
          reg681 = $signed($signed(reg17));
        end
    end
  always
    @(posedge clk) begin
      reg682 = {reg43, reg56};
    end
  always
    @(posedge clk) begin
      reg683 <= reg11;
      reg684 = reg17[(1'h0):(1'h0)];
      reg685 = (({(reg684[(1'h1):(1'h1)] >= wire4[(4'ha):(1'h1)])} ?
              (^~(+(!reg34))) : {(8'hb1), (&reg6)}) ?
          reg6[(5'h10):(4'he)] : wire2[(2'h2):(2'h2)]);
      reg686 = ({$unsigned($signed((-reg52)))} + $signed(wire4[(4'ha):(3'h5)]));
    end
  always
    @(posedge clk) begin
      reg687 <= wire70[(1'h1):(1'h0)];
      reg688 = (reg30[(1'h0):(1'h0)] + $signed((~&{reg55,
          (reg42 ? reg11 : reg69)})));
      reg689 <= (-(~(8'hb1)));
    end
  assign wire690 = {reg689[(2'h3):(1'h1)]};
  assign wire691 = (-(((|(reg65 ? reg56 : reg51)) | reg34) ?
                       reg6[(3'h5):(2'h3)] : (|{reg15})));
  always
    @(posedge clk) begin
      for (forvar692 = (1'h0); (forvar692 < (3'h4)); forvar692 = (forvar692 + (1'h1)))
        begin
          reg693 <= reg24;
          reg694 <= (+(~$unsigned((!(reg687 || wire2)))));
          reg695 = ((&(!(((8'hb8) ?
              reg36 : wire670) < (wire690 ^ wire670)))) ^ $unsigned(wire691[(2'h2):(1'h1)]));
          for (forvar696 = (1'h0); (forvar696 < (1'h1)); forvar696 = (forvar696 + (1'h1)))
            begin
              reg697 <= $signed($unsigned(reg23));
              reg698 <= (~&(-(reg10[(1'h0):(1'h0)] ?
                  (reg672 != (reg6 ?
                      reg54 : wire4)) : $signed($unsigned(wire691)))));
              reg699 <= ((~((!reg29) | wire2)) ?
                  $signed(forvar692) : reg49[(3'h4):(2'h2)]);
              reg700 = $signed((({(+reg694),
                  (8'hb7)} & reg18[(1'h1):(1'h0)]) | ($unsigned((wire4 ?
                  reg66 : reg56)) >> $signed((forvar696 ? reg57 : reg29)))));
            end
          reg701 <= $unsigned($signed($signed((reg31 <<< (reg12 ?
              (8'h9d) : reg6)))));
        end
      reg702 <= (~^reg43[(4'hf):(3'h7)]);
      if ((+{reg694, $signed((((8'h9d) <= wire71) - reg702[(3'h6):(3'h4)]))}))
        begin
          reg703 = $signed(reg19);
        end
      else
        begin
          reg704 <= reg61;
        end
      reg705 = $unsigned({reg689[(2'h3):(1'h0)], reg672});
      reg706 = (~|$signed(($signed((reg30 ?
          (7'h43) : reg15)) == reg65[(2'h2):(1'h0)])));
    end
  always
    @(posedge clk) begin
      if ($unsigned($unsigned(reg52[(1'h0):(1'h0)])))
        begin
          reg707 <= reg42;
        end
      else
        begin
          reg707 <= (~&(({$signed(reg17), (reg702 ? reg683 : reg687)} ?
                  $signed({wire70, (8'hb8)}) : (!(reg69 ? reg43 : reg15))) ?
              (((8'hab) || $signed(reg693)) ?
                  $unsigned(reg676[(2'h2):(1'h0)]) : reg22) : $unsigned($signed(reg49))));
          reg708 <= $unsigned(reg31);
        end
      reg709 <= ($unsigned(reg69) ?
          $unsigned({$signed($unsigned(reg22)),
              $signed((~^reg701))}) : {($unsigned({wire4, reg687}) ?
                  (~&wire1[(3'h4):(1'h1)]) : ((wire691 ^ reg42) ?
                      wire2[(2'h2):(1'h1)] : $signed(reg702)))});
      for (forvar710 = (1'h0); (forvar710 < (3'h4)); forvar710 = (forvar710 + (1'h1)))
        begin
          reg711 <= (reg39 ?
              (reg701[(1'h1):(1'h0)] ?
                  (reg702 ?
                      reg69 : $signed(reg19[(1'h1):(1'h1)])) : (~|reg708)) : ($signed($unsigned($signed(reg708))) >>> (&((~|reg61) ^ $signed((8'hb3))))));
          reg712 = $signed($signed({$signed((|reg56))}));
          reg713 <= {(8'ha3), $unsigned({$signed((reg6 ? reg8 : reg66))})};
          for (forvar714 = (1'h0); (forvar714 < (1'h0)); forvar714 = (forvar714 + (1'h1)))
            begin
              reg715 = reg56;
              reg716 = wire1[(4'hc):(4'h8)];
              reg717 = {($unsigned(reg29[(2'h2):(1'h0)]) ?
                      $unsigned($signed(reg12[(1'h0):(1'h0)])) : (8'hac))};
              reg718 <= (-($unsigned(({reg24, (8'hba)} ? {reg23} : reg34)) ?
                  $signed(reg63) : reg19));
              reg719 <= reg713;
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module463
#(parameter param669 = ((((((8'ha6) ? (8'hb2) : (8'hb8)) - {(8'ha1)}) ? (((8'hb5) ? (8'hab) : (8'ha1)) >>> ((7'h42) < (8'hb1))) : {{(7'h43)}, (|(8'hb8))}) ? (~&(((8'hb5) || (8'ha6)) && ((8'hbb) + (8'hbe)))) : (((8'ha0) ? ((8'ha2) ? (8'haf) : (8'hb4)) : ((8'h9f) ? (8'hb5) : (8'hab))) ? (((8'hb7) ? (7'h41) : (8'hbf)) <= ((8'hb6) ? (8'hba) : (8'ha3))) : {((8'ha1) ? (8'h9d) : (8'ha5))})) ? ((~|((&(8'hb5)) ? ((8'hbf) && (8'ha9)) : ((8'hae) | (8'ha9)))) | ((((8'ha0) ? (8'hb6) : (8'haf)) ? ((8'hbd) ? (8'hb8) : (8'hb0)) : (+(8'ha0))) ? {(!(8'ha3))} : (((8'haf) * (8'hac)) ? {(8'had)} : (~^(8'hb8))))) : (+{(|(|(8'haf)))})))
(y, clk, wire467, wire466, wire465, wire464);
  output wire [(32'h90c):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(4'hd):(1'h0)] wire467;
  input wire signed [(5'h15):(1'h0)] wire466;
  input wire signed [(2'h2):(1'h0)] wire465;
  input wire [(4'hd):(1'h0)] wire464;
  wire [(5'h11):(1'h0)] wire547;
  wire [(5'h10):(1'h0)] wire471;
  reg [(2'h2):(1'h0)] reg668 = (1'h0);
  reg [(3'h7):(1'h0)] reg667 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg666 = (1'h0);
  reg [(3'h6):(1'h0)] reg665 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg662 = (1'h0);
  reg [(5'h10):(1'h0)] reg660 = (1'h0);
  reg [(4'h8):(1'h0)] reg658 = (1'h0);
  reg [(5'h15):(1'h0)] reg657 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg653 = (1'h0);
  reg [(2'h2):(1'h0)] reg650 = (1'h0);
  reg [(4'hc):(1'h0)] reg649 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg648 = (1'h0);
  reg [(4'hd):(1'h0)] reg645 = (1'h0);
  reg [(3'h5):(1'h0)] reg643 = (1'h0);
  reg [(3'h6):(1'h0)] reg642 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg641 = (1'h0);
  reg [(4'ha):(1'h0)] reg629 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg627 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg626 = (1'h0);
  reg [(2'h2):(1'h0)] reg623 = (1'h0);
  reg [(5'h14):(1'h0)] reg622 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg621 = (1'h0);
  reg [(2'h3):(1'h0)] reg620 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg615 = (1'h0);
  reg [(4'hd):(1'h0)] reg613 = (1'h0);
  reg [(3'h5):(1'h0)] reg611 = (1'h0);
  reg [(4'h9):(1'h0)] reg608 = (1'h0);
  reg [(5'h14):(1'h0)] reg607 = (1'h0);
  reg [(4'ha):(1'h0)] reg606 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg605 = (1'h0);
  reg [(4'hb):(1'h0)] reg604 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg602 = (1'h0);
  reg [(4'hd):(1'h0)] reg600 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg599 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg597 = (1'h0);
  reg [(5'h10):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg593 = (1'h0);
  reg [(3'h4):(1'h0)] reg592 = (1'h0);
  reg [(2'h2):(1'h0)] reg585 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg583 = (1'h0);
  reg [(4'hd):(1'h0)] reg580 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg579 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg577 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg576 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg575 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg572 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg571 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg569 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg565 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg562 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg561 = (1'h0);
  reg [(5'h15):(1'h0)] reg560 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg559 = (1'h0);
  reg [(4'he):(1'h0)] reg556 = (1'h0);
  reg [(5'h10):(1'h0)] reg553 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg552 = (1'h0);
  reg [(5'h12):(1'h0)] reg551 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg549 = (1'h0);
  reg [(5'h10):(1'h0)] reg545 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg544 = (1'h0);
  reg [(2'h2):(1'h0)] reg543 = (1'h0);
  reg [(4'hf):(1'h0)] reg531 = (1'h0);
  reg [(4'hf):(1'h0)] reg530 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg527 = (1'h0);
  reg [(4'hb):(1'h0)] reg526 = (1'h0);
  reg [(4'he):(1'h0)] reg521 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg519 = (1'h0);
  reg [(2'h3):(1'h0)] reg518 = (1'h0);
  reg [(5'h12):(1'h0)] reg517 = (1'h0);
  reg [(4'hf):(1'h0)] reg515 = (1'h0);
  reg [(5'h15):(1'h0)] reg514 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg512 = (1'h0);
  reg [(3'h6):(1'h0)] reg510 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg508 = (1'h0);
  reg [(3'h5):(1'h0)] reg507 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg505 = (1'h0);
  reg [(5'h14):(1'h0)] reg504 = (1'h0);
  reg [(4'ha):(1'h0)] reg503 = (1'h0);
  reg [(4'hf):(1'h0)] reg502 = (1'h0);
  reg [(4'hf):(1'h0)] reg501 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg500 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg497 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg494 = (1'h0);
  reg [(4'hd):(1'h0)] reg491 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg488 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg487 = (1'h0);
  reg [(5'h15):(1'h0)] reg483 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg482 = (1'h0);
  reg [(2'h2):(1'h0)] reg481 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg478 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg477 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg476 = (1'h0);
  reg [(4'ha):(1'h0)] reg475 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg474 = (1'h0);
  reg [(4'h8):(1'h0)] reg470 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg468 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg664 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg663 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg661 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar659 = (1'h0);
  reg [(5'h12):(1'h0)] forvar656 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg655 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg654 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar645 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg652 = (1'h0);
  reg [(4'he):(1'h0)] reg651 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg647 = (1'h0);
  reg [(4'hf):(1'h0)] reg646 = (1'h0);
  reg [(3'h5):(1'h0)] reg644 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg640 = (1'h0);
  reg [(4'h9):(1'h0)] reg639 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg638 = (1'h0);
  reg [(4'he):(1'h0)] forvar637 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg636 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg635 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg634 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg633 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg632 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg631 = (1'h0);
  reg [(3'h6):(1'h0)] forvar630 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg628 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar625 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg624 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar619 = (1'h0);
  reg [(5'h13):(1'h0)] forvar618 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg617 = (1'h0);
  reg [(5'h15):(1'h0)] reg616 = (1'h0);
  reg signed [(4'he):(1'h0)] reg614 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg612 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar610 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg609 = (1'h0);
  reg [(3'h6):(1'h0)] forvar603 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg601 = (1'h0);
  reg [(2'h3):(1'h0)] forvar598 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg596 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar594 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg591 = (1'h0);
  reg [(5'h15):(1'h0)] forvar590 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg589 = (1'h0);
  reg [(4'h8):(1'h0)] forvar588 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg587 = (1'h0);
  reg [(4'hc):(1'h0)] reg586 = (1'h0);
  reg [(4'h8):(1'h0)] forvar584 = (1'h0);
  reg [(5'h11):(1'h0)] forvar582 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg581 = (1'h0);
  reg [(4'hf):(1'h0)] reg578 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar574 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg573 = (1'h0);
  reg [(3'h6):(1'h0)] reg570 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg568 = (1'h0);
  reg [(4'ha):(1'h0)] reg567 = (1'h0);
  reg [(2'h2):(1'h0)] forvar566 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar564 = (1'h0);
  reg [(5'h10):(1'h0)] reg563 = (1'h0);
  reg [(3'h6):(1'h0)] reg558 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg557 = (1'h0);
  reg [(5'h14):(1'h0)] forvar555 = (1'h0);
  reg [(3'h7):(1'h0)] forvar554 = (1'h0);
  reg [(4'hf):(1'h0)] reg550 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar548 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg546 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg542 = (1'h0);
  reg [(5'h13):(1'h0)] reg541 = (1'h0);
  reg [(3'h6):(1'h0)] forvar540 = (1'h0);
  reg [(4'hc):(1'h0)] reg539 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg538 = (1'h0);
  reg [(5'h10):(1'h0)] forvar537 = (1'h0);
  reg [(5'h11):(1'h0)] forvar536 = (1'h0);
  reg [(4'ha):(1'h0)] reg535 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg534 = (1'h0);
  reg [(4'hb):(1'h0)] reg533 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg532 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg529 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar528 = (1'h0);
  reg [(3'h6):(1'h0)] reg525 = (1'h0);
  reg [(4'hd):(1'h0)] reg524 = (1'h0);
  reg [(5'h15):(1'h0)] forvar523 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar522 = (1'h0);
  reg [(5'h15):(1'h0)] reg520 = (1'h0);
  reg [(5'h11):(1'h0)] reg516 = (1'h0);
  reg signed [(4'he):(1'h0)] reg513 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar511 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg506 = (1'h0);
  reg [(5'h10):(1'h0)] reg509 = (1'h0);
  reg [(4'h9):(1'h0)] forvar506 = (1'h0);
  reg signed [(4'he):(1'h0)] reg499 = (1'h0);
  reg [(3'h6):(1'h0)] reg498 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg496 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg495 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg493 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg492 = (1'h0);
  reg [(5'h12):(1'h0)] forvar490 = (1'h0);
  reg [(3'h6):(1'h0)] forvar489 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg486 = (1'h0);
  reg [(4'hf):(1'h0)] reg485 = (1'h0);
  reg [(3'h4):(1'h0)] forvar484 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg480 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg479 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg473 = (1'h0);
  reg [(4'hf):(1'h0)] forvar472 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg469 = (1'h0);
  assign y = {wire547,
                 wire471,
                 reg668,
                 reg667,
                 reg666,
                 reg665,
                 reg662,
                 reg660,
                 reg658,
                 reg657,
                 reg653,
                 reg650,
                 reg649,
                 reg648,
                 reg645,
                 reg643,
                 reg642,
                 reg641,
                 reg629,
                 reg627,
                 reg626,
                 reg623,
                 reg622,
                 reg621,
                 reg620,
                 reg615,
                 reg613,
                 reg611,
                 reg608,
                 reg607,
                 reg606,
                 reg605,
                 reg604,
                 reg602,
                 reg600,
                 reg599,
                 reg597,
                 reg595,
                 reg593,
                 reg592,
                 reg585,
                 reg583,
                 reg580,
                 reg579,
                 reg577,
                 reg576,
                 reg575,
                 reg572,
                 reg571,
                 reg569,
                 reg565,
                 reg562,
                 reg561,
                 reg560,
                 reg559,
                 reg556,
                 reg553,
                 reg552,
                 reg551,
                 reg549,
                 reg545,
                 reg544,
                 reg543,
                 reg531,
                 reg530,
                 reg527,
                 reg526,
                 reg521,
                 reg519,
                 reg518,
                 reg517,
                 reg515,
                 reg514,
                 reg512,
                 reg510,
                 reg508,
                 reg507,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 reg501,
                 reg500,
                 reg497,
                 reg494,
                 reg491,
                 reg488,
                 reg487,
                 reg483,
                 reg482,
                 reg481,
                 reg478,
                 reg477,
                 reg476,
                 reg475,
                 reg474,
                 reg470,
                 reg468,
                 reg664,
                 reg663,
                 reg661,
                 forvar659,
                 forvar656,
                 reg655,
                 reg654,
                 forvar645,
                 reg652,
                 reg651,
                 reg647,
                 reg646,
                 reg644,
                 reg640,
                 reg639,
                 reg638,
                 forvar637,
                 reg636,
                 reg635,
                 reg634,
                 reg633,
                 reg632,
                 reg631,
                 forvar630,
                 reg628,
                 forvar625,
                 reg624,
                 forvar619,
                 forvar618,
                 reg617,
                 reg616,
                 reg614,
                 reg612,
                 forvar610,
                 reg609,
                 forvar603,
                 reg601,
                 forvar598,
                 reg596,
                 forvar594,
                 reg591,
                 forvar590,
                 reg589,
                 forvar588,
                 reg587,
                 reg586,
                 forvar584,
                 forvar582,
                 reg581,
                 reg578,
                 forvar574,
                 reg573,
                 reg570,
                 reg568,
                 reg567,
                 forvar566,
                 forvar564,
                 reg563,
                 reg558,
                 reg557,
                 forvar555,
                 forvar554,
                 reg550,
                 forvar548,
                 reg546,
                 reg542,
                 reg541,
                 forvar540,
                 reg539,
                 reg538,
                 forvar537,
                 forvar536,
                 reg535,
                 reg534,
                 reg533,
                 reg532,
                 reg529,
                 forvar528,
                 reg525,
                 reg524,
                 forvar523,
                 forvar522,
                 reg520,
                 reg516,
                 reg513,
                 forvar511,
                 reg506,
                 reg509,
                 forvar506,
                 reg499,
                 reg498,
                 reg496,
                 reg495,
                 reg493,
                 reg492,
                 forvar490,
                 forvar489,
                 reg486,
                 reg485,
                 forvar484,
                 reg480,
                 reg479,
                 reg473,
                 forvar472,
                 reg469,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg468 <= wire467[(2'h2):(1'h0)];
      reg469 = wire467[(1'h0):(1'h0)];
      reg470 <= (8'ha4);
    end
  assign wire471 = reg468[(3'h4):(2'h2)];
  always
    @(posedge clk) begin
      for (forvar472 = (1'h0); (forvar472 < (2'h2)); forvar472 = (forvar472 + (1'h1)))
        begin
          reg473 = reg470[(3'h6):(1'h0)];
          reg474 <= {(wire465 >> wire466),
              ((wire471 ?
                  $unsigned({reg468}) : ((reg473 ? wire465 : wire465) ?
                      $signed(wire467) : (wire464 & wire464))) && wire464)};
          reg475 <= ($signed(reg473) * reg468[(1'h1):(1'h0)]);
          if (({wire466[(5'h15):(5'h10)],
              $signed($signed(wire466[(1'h1):(1'h0)]))} != wire465[(1'h0):(1'h0)]))
            begin
              reg476 <= wire471[(3'h6):(3'h6)];
              reg477 <= $signed((8'ha0));
              reg478 <= reg474;
              reg479 = (~&($signed($signed((reg474 ^ reg478))) && ($signed($unsigned((8'hbf))) <<< (forvar472 - $signed(reg475)))));
            end
          else
            begin
              reg479 = (~^({$unsigned((^reg474)),
                  $unsigned(((7'h42) ?
                      reg474 : reg478))} > $signed(reg470[(3'h7):(2'h3)])));
              reg480 = {($signed(({wire465} + reg474[(3'h4):(2'h3)])) ?
                      wire471[(4'h9):(3'h6)] : (wire471[(5'h10):(3'h4)] < forvar472))};
              reg481 <= (|(^~$unsigned(((8'h9c) == (8'ha8)))));
              reg482 <= $unsigned({reg480[(2'h2):(1'h1)]});
              reg483 <= reg468;
            end
          for (forvar484 = (1'h0); (forvar484 < (1'h0)); forvar484 = (forvar484 + (1'h1)))
            begin
              reg485 = ((|$signed($unsigned((wire466 ~^ wire467)))) & (reg476 ~^ $unsigned((forvar472[(4'hf):(4'hf)] ?
                  reg481 : $signed(forvar472)))));
              reg486 = reg475[(3'h7):(3'h7)];
            end
        end
      reg487 <= (+{$signed({(&reg483), (reg473 ? wire465 : reg481)})});
      reg488 <= reg477;
      for (forvar489 = (1'h0); (forvar489 < (2'h2)); forvar489 = (forvar489 + (1'h1)))
        begin
          for (forvar490 = (1'h0); (forvar490 < (2'h2)); forvar490 = (forvar490 + (1'h1)))
            begin
              reg491 <= ((~&{(8'hb5),
                  $signed((reg474 ?
                      reg480 : reg468))}) + ($unsigned($signed((reg474 ?
                  reg479 : reg486))) >= (wire466[(4'hf):(3'h5)] > {wire464[(4'hc):(2'h3)],
                  $signed(forvar489)})));
              reg492 = (forvar484[(2'h3):(1'h0)] ^~ ((reg481 & (~&(forvar489 + reg468))) ?
                  $unsigned($signed(forvar489)) : (($unsigned(reg476) >>> $unsigned(forvar472)) + reg481[(1'h0):(1'h0)])));
              reg493 = reg485;
              reg494 <= $unsigned((forvar484 + (reg470 ^~ (forvar484[(1'h0):(1'h0)] ?
                  (reg481 << reg479) : (wire471 ? reg486 : reg474)))));
            end
          if ((&$signed(reg487[(4'hb):(3'h7)])))
            begin
              reg495 = reg493;
              reg496 = reg491;
              reg497 <= (((($unsigned(wire465) ?
                      {forvar484,
                          forvar489} : reg482) <<< {reg480[(4'hc):(1'h1)]}) ?
                  reg476[(4'h9):(4'h9)] : $signed((~&reg495))) == ($unsigned(({reg480,
                      wire471} & $signed(reg493))) ?
                  {(wire464[(1'h1):(1'h1)] | $unsigned((8'hac)))} : (!reg476[(2'h3):(2'h2)])));
              reg498 = $signed(reg468);
            end
          else
            begin
              reg497 <= {(~$signed($unsigned(wire466[(5'h10):(4'ha)])))};
              reg498 = $signed($unsigned((~reg498[(3'h4):(2'h2)])));
              reg499 = $unsigned($unsigned(($unsigned($signed(reg476)) | $unsigned($signed((8'ha6))))));
              reg500 <= (-$unsigned((reg487[(4'h9):(1'h0)] >> (reg468[(3'h7):(3'h6)] <<< {reg497}))));
              reg501 <= ((^~reg482[(2'h2):(2'h2)]) == $unsigned(forvar484));
            end
          if ((reg492 > (|($unsigned((reg494 - (8'hb1))) <= (reg479 ?
              reg501[(4'hc):(3'h4)] : $signed(reg499))))))
            begin
              reg502 <= $unsigned(($signed(reg483) ?
                  $signed(reg491) : {((reg481 ^ reg475) * $signed(reg468)),
                      $unsigned($unsigned(reg479))}));
              reg503 <= $unsigned((~^($signed($unsigned(reg475)) ?
                  $signed($unsigned(reg487)) : ((7'h42) | ((7'h40) ?
                      reg492 : forvar472)))));
              reg504 <= (7'h42);
              reg505 <= (($unsigned(reg479) ?
                  $signed(reg468) : $signed(($signed(reg491) > ((8'ha2) ?
                      reg480 : reg477)))) >= $signed(((~^(&reg499)) ?
                  reg473[(2'h3):(1'h0)] : (8'ha9))));
            end
          else
            begin
              reg502 <= $signed({$signed((~|reg483))});
              reg503 <= $signed($signed((reg477[(4'hd):(4'hc)] ?
                  ((reg492 - reg485) ? reg492 : $unsigned(reg475)) : ({reg480} ?
                      $unsigned(reg501) : forvar472))));
              reg504 <= ($signed(reg491[(1'h1):(1'h0)]) ?
                  $unsigned((((^~(8'ha3)) ?
                      (reg481 < reg485) : ((8'hb5) == reg482)) || reg502)) : ($signed((wire464 ?
                      (8'h9e) : reg501)) >> $unsigned(reg483[(2'h2):(1'h0)])));
              reg505 <= (&(($signed(wire471) && ($signed((8'hab)) <= $signed(reg500))) ?
                  {wire466[(4'h8):(3'h7)]} : (((wire471 <= (8'ha8)) * $signed(reg482)) ?
                      $unsigned(reg500) : ((reg496 < (8'hbb)) == reg470))));
            end
        end
    end
  always
    @(posedge clk) begin
      if (($signed((reg468[(1'h1):(1'h0)] ?
          {{reg475, reg482}} : ((reg502 && wire464) ?
              $signed(reg478) : ((7'h40) && reg501)))) >> (~&wire471[(5'h10):(5'h10)])))
        begin
          for (forvar506 = (1'h0); (forvar506 < (2'h2)); forvar506 = (forvar506 + (1'h1)))
            begin
              reg507 <= (reg488 ?
                  ($unsigned($signed((wire467 ? wire467 : (8'ha6)))) ?
                      reg504[(3'h5):(1'h0)] : {(~&(reg474 ^~ reg505)),
                          ((reg500 ? wire465 : reg482) ?
                              (^wire467) : (~^reg468))}) : $unsigned(reg501[(4'h9):(4'h9)]));
              reg508 <= $signed(((($unsigned(reg474) ?
                      reg474[(4'hf):(4'h8)] : wire471) ?
                  $signed(reg474[(4'hf):(4'he)]) : (8'h9f)) > {reg475[(2'h2):(2'h2)],
                  ((8'hac) ? $signed(wire467) : (wire465 ? reg475 : reg494))}));
              reg509 = ((^~(~&{{reg483}})) & reg468);
            end
          reg510 <= ($unsigned({wire464[(4'ha):(4'h8)]}) == $signed(reg477[(2'h3):(2'h3)]));
        end
      else
        begin
          if ($signed(reg502[(4'h9):(2'h2)]))
            begin
              reg506 = $unsigned($signed((~|(^(8'hb3)))));
              reg507 <= ({(!$unsigned($unsigned(wire464))),
                      reg477[(5'h10):(4'h9)]} ?
                  (($unsigned((reg494 ^~ reg502)) ?
                          (reg505[(1'h0):(1'h0)] ^~ $signed(reg507)) : ($unsigned(wire471) & $signed(reg476))) ?
                      wire466 : $unsigned($unsigned((reg477 >> reg474)))) : (|($unsigned(reg478) ?
                      $signed($signed(reg470)) : ((-reg470) >> $signed(reg488)))));
              reg508 <= {(reg505[(3'h6):(1'h1)] >>> reg474[(4'ha):(3'h5)]),
                  $unsigned(reg474)};
            end
          else
            begin
              reg507 <= reg483[(1'h0):(1'h0)];
            end
          reg510 <= (wire467[(3'h4):(2'h3)] > (~reg488[(3'h4):(1'h1)]));
          for (forvar511 = (1'h0); (forvar511 < (1'h0)); forvar511 = (forvar511 + (1'h1)))
            begin
              reg512 <= reg500;
              reg513 = reg502;
              reg514 <= $signed($unsigned((^~$unsigned(((8'ha1) ?
                  (8'had) : reg506)))));
            end
        end
      reg515 <= $unsigned({$signed($unsigned(reg502[(4'h8):(1'h0)])),
          (-reg502)});
      reg516 = ((~^$unsigned(reg494[(1'h1):(1'h0)])) ?
          (((((8'hb5) ? reg500 : (8'ha3)) ?
                  (reg514 ? reg505 : reg494) : (reg478 ?
                      reg500 : wire466)) < reg500[(3'h5):(3'h5)]) ?
              (^~(~reg476)) : $unsigned($unsigned({reg483}))) : {($unsigned($signed(reg515)) ?
                  reg475[(4'ha):(3'h6)] : reg515[(4'hc):(4'h8)])});
      reg517 <= $signed(reg488[(4'ha):(3'h6)]);
    end
  always
    @(posedge clk) begin
      reg518 <= $unsigned($unsigned($signed(reg507[(3'h4):(2'h3)])));
      if (reg478[(2'h3):(2'h3)])
        begin
          reg519 <= {(reg481 ?
                  (($unsigned(reg504) >>> (reg508 ?
                      (8'hb3) : reg468)) || ((reg481 <<< reg504) ?
                      $unsigned(reg470) : reg501)) : reg501),
              (({reg507} <= ($unsigned(reg515) ?
                  reg515[(1'h0):(1'h0)] : $unsigned(wire471))) >> (!{(wire465 - reg470),
                  (^reg483)}))};
          reg520 = $unsigned(($signed(wire471[(3'h6):(2'h3)]) <= {($signed(reg468) == ((8'hac) | reg468)),
              $signed(reg515[(3'h4):(1'h0)])}));
          reg521 <= (~^reg483[(3'h7):(1'h0)]);
        end
      else
        begin
          reg520 = (wire465 ?
              ({(reg468 || reg474)} ?
                  $signed((reg481[(1'h1):(1'h1)] ?
                      (~reg497) : (|reg470))) : (((&reg478) <= reg512[(4'he):(3'h7)]) * reg477[(1'h1):(1'h1)])) : (reg487[(4'h8):(4'h8)] <= ((+$unsigned(reg468)) ^ ($unsigned(reg517) ?
                  $signed((7'h43)) : (-wire466)))));
        end
      for (forvar522 = (1'h0); (forvar522 < (2'h3)); forvar522 = (forvar522 + (1'h1)))
        begin
          for (forvar523 = (1'h0); (forvar523 < (1'h0)); forvar523 = (forvar523 + (1'h1)))
            begin
              reg524 = ((({$unsigned((8'hb7))} & $unsigned((wire465 ?
                  reg504 : (8'ha8)))) * reg510) ^~ $unsigned($signed(reg483)));
              reg525 = (~((|wire465[(2'h2):(1'h1)]) ?
                  ((~&(|wire466)) <<< wire464) : reg518));
              reg526 <= reg491;
              reg527 <= reg517[(2'h2):(1'h0)];
            end
          for (forvar528 = (1'h0); (forvar528 < (3'h4)); forvar528 = (forvar528 + (1'h1)))
            begin
              reg529 = (wire466[(2'h3):(2'h3)] < {((|reg478) ?
                      (^reg521) : ((reg521 ?
                          reg518 : reg488) << (reg470 | reg470)))});
            end
          if (wire471[(3'h7):(3'h5)])
            begin
              reg530 <= $unsigned($unsigned(($signed((!reg529)) != (^~$unsigned(reg497)))));
              reg531 <= wire464;
              reg532 = reg504;
            end
          else
            begin
              reg530 <= $unsigned(((($signed(reg532) << reg501[(3'h6):(2'h3)]) ?
                  ({reg504} ?
                      (forvar528 <= wire465) : (reg502 ?
                          reg504 : reg518)) : reg470) >= ((reg515 ?
                      {reg527} : (~|reg532)) ?
                  $unsigned((|reg494)) : $unsigned({reg529, reg483}))));
            end
          reg533 = (($signed(((+reg512) ^ ((7'h44) <<< reg474))) ~^ ((^{reg508,
                  reg520}) ?
              (~&(+wire466)) : $unsigned((reg527 - reg515)))) < $signed(forvar522));
          reg534 = {{$unsigned($signed(((8'h9d) ? reg500 : reg502)))}, reg476};
        end
      reg535 = reg530[(3'h5):(2'h2)];
    end
  always
    @(posedge clk) begin
      for (forvar536 = (1'h0); (forvar536 < (1'h1)); forvar536 = (forvar536 + (1'h1)))
        begin
          for (forvar537 = (1'h0); (forvar537 < (1'h0)); forvar537 = (forvar537 + (1'h1)))
            begin
              reg538 = (!reg487);
              reg539 = $unsigned({(reg488 ?
                      reg508[(3'h7):(1'h0)] : $signed($signed(reg512)))});
            end
          for (forvar540 = (1'h0); (forvar540 < (1'h0)); forvar540 = (forvar540 + (1'h1)))
            begin
              reg541 = $signed((~&({{reg514, reg470},
                  $unsigned(reg521)} < {((8'hb5) && reg491),
                  ((8'hb9) ? forvar537 : forvar540)})));
              reg542 = reg507;
              reg543 <= reg488;
              reg544 <= $signed($unsigned(reg491));
            end
        end
      reg545 <= ($unsigned(({{forvar537, reg500}, (&(8'hbe))} ?
          (^$unsigned(reg491)) : ($signed(reg544) ?
              (~&forvar537) : reg518[(2'h3):(2'h3)]))) <= reg542);
      reg546 = ($unsigned($signed(reg468)) <= reg494[(1'h1):(1'h0)]);
    end
  assign wire547 = $unsigned(reg468);
  always
    @(posedge clk) begin
      for (forvar548 = (1'h0); (forvar548 < (2'h3)); forvar548 = (forvar548 + (1'h1)))
        begin
          reg549 <= ((!(^$signed((~^reg510)))) ?
              (|($unsigned((reg517 >> reg475)) * $unsigned($unsigned(reg501)))) : ((+$signed(reg502)) ?
                  (reg544[(4'hb):(4'h8)] ?
                      $unsigned($unsigned(reg488)) : (~&reg510[(3'h5):(2'h3)])) : forvar548));
          reg550 = (|reg491[(4'ha):(1'h1)]);
          reg551 <= $unsigned(({(reg517 == (+reg544))} < $unsigned({reg512[(4'hc):(4'h8)]})));
          reg552 <= reg510;
          reg553 <= reg505[(3'h6):(3'h4)];
        end
      for (forvar554 = (1'h0); (forvar554 < (1'h0)); forvar554 = (forvar554 + (1'h1)))
        begin
          for (forvar555 = (1'h0); (forvar555 < (1'h0)); forvar555 = (forvar555 + (1'h1)))
            begin
              reg556 <= $unsigned(reg530);
              reg557 = $signed($unsigned($signed(wire466[(1'h1):(1'h0)])));
              reg558 = (-reg508);
              reg559 <= (~&(^{({reg508} <<< (reg497 ? reg507 : reg518)),
                  reg519[(4'ha):(3'h7)]}));
            end
          reg560 <= (~reg470);
          reg561 <= reg526[(2'h2):(2'h2)];
          reg562 <= reg557;
        end
      reg563 = (|$signed({(~|reg475)}));
      for (forvar564 = (1'h0); (forvar564 < (1'h0)); forvar564 = (forvar564 + (1'h1)))
        begin
          reg565 <= {reg527};
          for (forvar566 = (1'h0); (forvar566 < (2'h3)); forvar566 = (forvar566 + (1'h1)))
            begin
              reg567 = $unsigned($signed((reg517 ^~ ((reg551 ?
                      reg545 : forvar554) ?
                  (!reg470) : $unsigned(wire467)))));
              reg568 = (((!{(^~reg468), (^reg526)}) ?
                      {(7'h44)} : ({wire464[(4'hd):(3'h6)],
                              $unsigned((7'h40))} ?
                          {reg470[(1'h1):(1'h1)]} : {(wire547 >> reg482),
                              (-reg567)})) ?
                  $signed(reg501[(4'hb):(1'h0)]) : (8'hbe));
              reg569 <= (reg502[(3'h7):(2'h3)] <<< (~&((reg487 & reg508) ^ $signed((&reg470)))));
              reg570 = ((reg565[(3'h6):(3'h4)] ^ $signed(reg556[(1'h1):(1'h0)])) ?
                  ($unsigned($unsigned((&reg483))) && ($unsigned($unsigned(wire471)) ?
                      ($signed((8'hbe)) == reg508[(2'h2):(1'h1)]) : (~(reg518 * reg557)))) : $unsigned((+$signed((+reg508)))));
              reg571 <= (^~$signed($unsigned((reg468 < (reg544 ?
                  reg491 : (8'hb1))))));
            end
          reg572 <= (^(~reg503[(4'h9):(3'h4)]));
          reg573 = ($unsigned($signed(((reg481 - (8'hb7)) >>> (reg571 - reg527)))) <<< (((~^(+wire467)) >>> ($unsigned((8'ha8)) > $unsigned(forvar555))) || reg526[(1'h1):(1'h0)]));
          for (forvar574 = (1'h0); (forvar574 < (1'h0)); forvar574 = (forvar574 + (1'h1)))
            begin
              reg575 <= $signed($unsigned($unsigned(reg482[(1'h1):(1'h0)])));
              reg576 <= (8'ha9);
              reg577 <= ((8'ha8) & (-reg507));
            end
        end
    end
  always
    @(posedge clk) begin
      reg578 = $signed($unsigned(($signed((reg515 ?
          reg527 : reg502)) >>> $signed((wire465 ~^ reg549)))));
      reg579 <= (-$unsigned(((|(wire471 ? (8'hb7) : reg510)) ?
          ($unsigned((7'h41)) ?
              reg562 : reg475[(2'h3):(2'h3)]) : (~^(reg517 ^~ reg512)))));
      reg580 <= reg503[(3'h6):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg581 = reg560[(5'h12):(4'hf)];
      for (forvar582 = (1'h0); (forvar582 < (1'h0)); forvar582 = (forvar582 + (1'h1)))
        begin
          reg583 <= $unsigned($unsigned($unsigned(reg556[(1'h0):(1'h0)])));
          for (forvar584 = (1'h0); (forvar584 < (3'h4)); forvar584 = (forvar584 + (1'h1)))
            begin
              reg585 <= $unsigned($unsigned($signed($signed((reg491 ?
                  reg491 : (8'ha2))))));
              reg586 = (-$unsigned({((reg491 ? reg530 : reg487) ?
                      (reg487 ? reg571 : reg549) : (reg577 ? reg510 : reg510)),
                  reg531[(4'hb):(2'h3)]}));
            end
          reg587 = {reg549[(2'h2):(1'h1)],
              (+$signed($signed(reg580[(2'h3):(2'h3)])))};
          for (forvar588 = (1'h0); (forvar588 < (2'h2)); forvar588 = (forvar588 + (1'h1)))
            begin
              reg589 = (^{($unsigned(reg587[(4'ha):(3'h5)]) ?
                      reg475[(2'h3):(1'h1)] : $signed($signed(reg507))),
                  (|$unsigned(reg559[(2'h3):(1'h1)]))});
            end
          for (forvar590 = (1'h0); (forvar590 < (3'h4)); forvar590 = (forvar590 + (1'h1)))
            begin
              reg591 = {($signed(($unsigned(wire471) > $unsigned(reg585))) ?
                      (8'ha4) : ($unsigned(reg531) ?
                          $unsigned((8'hb1)) : (^(reg530 ? reg561 : reg576)))),
                  (~(^reg474[(4'ha):(4'h8)]))};
              reg592 <= ($signed(reg556[(3'h7):(2'h3)]) * ($signed({(reg544 ?
                          reg586 : reg553),
                      $unsigned(reg526)}) ?
                  (reg521[(3'h7):(3'h7)] ?
                      $signed($signed(reg519)) : {$unsigned((7'h40))}) : reg530[(3'h6):(3'h4)]));
              reg593 <= ($unsigned($unsigned(reg545)) ?
                  (^reg507) : {($signed((&reg508)) && $unsigned($unsigned(reg507)))});
            end
        end
      for (forvar594 = (1'h0); (forvar594 < (1'h1)); forvar594 = (forvar594 + (1'h1)))
        begin
          reg595 <= $signed(reg515);
        end
    end
  always
    @(posedge clk) begin
      reg596 = ((reg497[(4'hb):(3'h6)] ?
              (($signed(reg515) >> (reg595 ?
                  reg488 : reg561)) > reg551[(3'h6):(3'h4)]) : {{reg569[(5'h15):(2'h2)],
                      reg477}}) ?
          reg507[(1'h0):(1'h0)] : {$signed($unsigned(reg501)),
              reg474[(4'h8):(1'h0)]});
      reg597 <= reg501[(1'h0):(1'h0)];
    end
  always
    @(posedge clk) begin
      for (forvar598 = (1'h0); (forvar598 < (2'h3)); forvar598 = (forvar598 + (1'h1)))
        begin
          if ({{$signed({(reg530 > reg545), (+reg507)}),
                  (^~(reg585[(2'h2):(2'h2)] ?
                      $signed(reg482) : $signed(reg474)))},
              reg494[(1'h1):(1'h1)]})
            begin
              reg599 <= ((8'hb8) ?
                  (reg565[(3'h5):(1'h0)] ?
                      $unsigned({reg572}) : $unsigned((reg497 ?
                          (reg531 ?
                              reg468 : reg478) : reg552[(1'h1):(1'h1)]))) : (forvar598[(1'h1):(1'h1)] < reg478[(1'h1):(1'h1)]));
              reg600 <= (~^(~^(($unsigned(reg544) <<< (reg530 >= reg545)) * (^(~|reg551)))));
              reg601 = (~^reg597[(1'h0):(1'h0)]);
              reg602 <= reg517;
            end
          else
            begin
              reg601 = ($signed(reg521[(4'hd):(4'hc)]) ?
                  (reg543[(1'h0):(1'h0)] ?
                      (|((reg572 ? reg477 : wire547) ?
                          (reg545 ? (8'ha7) : reg560) : reg559)) : (wire467 ?
                          {(^forvar598)} : $signed((|reg501)))) : (-(+reg600[(4'hb):(1'h1)])));
            end
          for (forvar603 = (1'h0); (forvar603 < (3'h4)); forvar603 = (forvar603 + (1'h1)))
            begin
              reg604 <= reg503[(1'h1):(1'h0)];
              reg605 <= $signed(($signed((~&(reg593 << reg579))) | $unsigned(reg514)));
              reg606 <= {$signed(reg507), reg601};
              reg607 <= reg517;
            end
          reg608 <= (~&($unsigned(reg501[(1'h0):(1'h0)]) | (+reg500[(2'h3):(1'h0)])));
          reg609 = $unsigned(($unsigned({(+reg530)}) != (~|$unsigned((8'hb5)))));
          for (forvar610 = (1'h0); (forvar610 < (3'h4)); forvar610 = (forvar610 + (1'h1)))
            begin
              reg611 <= (^~(reg576 ?
                  (^~$unsigned((reg531 <= reg543))) : $signed({{reg527},
                      (reg482 >= reg510)})));
              reg612 = reg501[(4'h8):(3'h6)];
              reg613 <= reg515;
              reg614 = (!$signed($unsigned(reg500[(1'h0):(1'h0)])));
              reg615 <= {reg575,
                  $signed({reg477,
                      ($unsigned(reg552) ?
                          (reg593 || wire465) : reg607[(3'h7):(3'h5)])})};
            end
        end
      reg616 = $unsigned($signed(forvar598));
      reg617 = wire467;
      for (forvar618 = (1'h0); (forvar618 < (1'h0)); forvar618 = (forvar618 + (1'h1)))
        begin
          for (forvar619 = (1'h0); (forvar619 < (1'h1)); forvar619 = (forvar619 + (1'h1)))
            begin
              reg620 <= (~&reg482);
              reg621 <= $signed((+(7'h43)));
              reg622 <= $unsigned(reg488[(3'h4):(2'h3)]);
              reg623 <= ({(~|forvar619[(3'h4):(3'h4)])} & (reg556 ?
                  $signed($signed($signed(reg600))) : {((^~reg585) ?
                          $unsigned(forvar598) : (reg549 ? reg617 : reg577))}));
              reg624 = ($signed((~((reg605 ? forvar603 : reg505) * reg494))) ?
                  $signed($signed($signed(reg477[(3'h4):(1'h1)]))) : ({((&reg526) > $signed(reg580)),
                      reg612} <= reg481));
            end
          for (forvar625 = (1'h0); (forvar625 < (1'h0)); forvar625 = (forvar625 + (1'h1)))
            begin
              reg626 <= (-(~&$unsigned(($signed(reg569) + reg543))));
              reg627 <= ($signed((reg497 ?
                  (-reg608[(2'h2):(1'h0)]) : $signed($unsigned(reg518)))) ^ (reg518[(2'h2):(1'h0)] + (8'hb2)));
              reg628 = reg622[(5'h13):(3'h5)];
              reg629 <= ($unsigned(((&reg614) ?
                  $signed($signed(reg628)) : (reg614[(4'ha):(3'h4)] ?
                      (reg561 - reg545) : reg620))) >= ({($signed(reg545) << (reg575 || reg481)),
                  (^reg561[(3'h4):(2'h2)])} >> $signed(({reg614,
                  reg622} ^ {reg577}))));
            end
          for (forvar630 = (1'h0); (forvar630 < (2'h3)); forvar630 = (forvar630 + (1'h1)))
            begin
              reg631 = ($unsigned($signed(({(8'haa), reg475} ?
                  ((8'ha6) ? (8'ha3) : reg616) : ((8'ha7) ?
                      (8'h9c) : forvar603)))) && ((|((reg549 ?
                          reg599 : wire467) ?
                      (reg514 ? reg549 : wire465) : (reg565 * reg577))) ?
                  $unsigned(reg477) : reg491[(1'h0):(1'h0)]));
              reg632 = ({(8'hbc), reg514[(4'h9):(1'h0)]} ?
                  (8'hab) : {(8'hb8), $unsigned($unsigned($signed((8'hb7))))});
              reg633 = reg593;
              reg634 = {$signed(($signed({wire466}) + (reg475 ^~ (+(8'hab)))))};
              reg635 = reg576[(4'h9):(2'h3)];
            end
          reg636 = ($signed((~&$signed(reg627))) ?
              (reg580 ?
                  $unsigned({$unsigned(reg572),
                      (reg616 ?
                          (8'hbd) : reg468)}) : $unsigned({reg614[(4'h8):(2'h2)],
                      reg620[(2'h3):(1'h0)]})) : (!reg607));
          for (forvar637 = (1'h0); (forvar637 < (3'h4)); forvar637 = (forvar637 + (1'h1)))
            begin
              reg638 = reg576;
              reg639 = reg604;
            end
        end
      reg640 = (^(^~((reg572 ? (^reg475) : (8'ha4)) ?
          reg527[(2'h2):(2'h2)] : ($signed(reg622) >= $unsigned(reg606)))));
    end
  always
    @(posedge clk) begin
      if (reg593[(4'hf):(2'h3)])
        begin
          reg641 <= (~(!$signed(((!reg606) ? (wire464 <<< reg597) : reg621))));
          if (($unsigned($signed(reg510)) >>> ($signed($unsigned((&(8'hb2)))) != ((reg544[(4'hf):(4'hb)] | $unsigned((8'hab))) ?
              (8'hac) : $unsigned(reg627)))))
            begin
              reg642 <= $unsigned($signed(($signed(reg605) << $unsigned((reg613 ?
                  reg602 : reg519)))));
              reg643 <= {({(reg476 || (^reg545))} + {(|$signed(reg531))}),
                  {reg597[(4'h9):(3'h7)]}};
              reg644 = (((((reg622 ? reg503 : reg517) >> (reg592 ?
                          wire547 : reg629)) ?
                      $unsigned((reg597 ?
                          (8'hbd) : reg530)) : (reg518[(2'h3):(1'h0)] << (8'had))) ?
                  reg569 : reg571) >> reg504);
            end
          else
            begin
              reg642 <= reg577[(3'h4):(2'h2)];
              reg644 = (~((~&((reg500 ?
                      reg500 : reg599) > (reg482 * (8'hb4)))) ?
                  $unsigned((reg510[(1'h1):(1'h1)] ^~ reg607[(5'h13):(4'h8)])) : ($signed(reg621) ?
                      reg615[(5'h12):(3'h4)] : {(!reg527)})));
              reg645 <= ($unsigned($signed({$unsigned((8'hb7))})) < ($signed($unsigned((^wire471))) ?
                  {{(reg599 & reg604),
                          (reg600 ?
                              reg512 : reg500)}} : $unsigned((~^(8'haf)))));
            end
          if (((reg583[(1'h0):(1'h0)] ?
                  $signed($unsigned(reg515[(3'h6):(2'h2)])) : reg605[(1'h0):(1'h0)]) ?
              {reg521[(1'h1):(1'h1)]} : (-((~&reg599[(5'h13):(3'h4)]) ?
                  ($signed(reg615) ?
                      reg482 : (reg481 ?
                          reg502 : reg642)) : (reg644[(2'h3):(1'h0)] <= $signed(reg622))))))
            begin
              reg646 = (reg491[(1'h1):(1'h0)] <= $unsigned(reg477));
              reg647 = $signed($signed(({$signed(reg505),
                  reg642} << reg474[(2'h3):(1'h0)])));
            end
          else
            begin
              reg648 <= reg643[(3'h5):(3'h5)];
              reg649 <= (&($signed((~&$unsigned(reg595))) ?
                  $signed((((8'hac) < reg487) ?
                      reg502 : $signed(reg579))) : wire471));
              reg650 <= reg527[(1'h1):(1'h0)];
              reg651 = {(^$unsigned(($unsigned(wire466) ?
                      {reg474, reg561} : (reg580 ? reg627 : reg552)))),
                  ($unsigned(($signed(reg606) ?
                      $unsigned(reg515) : (reg468 && reg608))) <= ({reg613[(4'hd):(2'h3)],
                      (wire464 ?
                          reg475 : reg650)} != ($signed(reg615) <= {reg497,
                      (8'ha5)})))};
            end
          reg652 = ((^~reg623) < reg565);
          reg653 <= $unsigned((((~reg623) ?
              {((8'hae) - reg580)} : ({reg604, reg478} ?
                  reg551[(1'h0):(1'h0)] : (reg475 ?
                      reg501 : reg512))) ^ (((-reg575) ?
                  reg559 : $signed((7'h41))) ?
              {$unsigned((8'hb9)), (&reg599)} : ({wire547} ?
                  (!(8'hb9)) : (reg599 ? reg559 : reg491)))));
        end
      else
        begin
          reg641 <= ($unsigned((((|(7'h43)) & {(8'hb3)}) ?
                  $unsigned(wire471) : reg527[(1'h1):(1'h0)])) ?
              reg608 : ({($signed((8'h9d)) < (&reg595)),
                      wire547[(4'hf):(1'h1)]} ?
                  reg607[(4'hd):(3'h7)] : $unsigned(reg500)));
          reg644 = $signed($unsigned({(~{(8'hb4)}),
              (reg650 ? reg652 : ((8'haa) ? reg543 : reg559))}));
          for (forvar645 = (1'h0); (forvar645 < (2'h3)); forvar645 = (forvar645 + (1'h1)))
            begin
              reg646 = $signed($signed(reg643));
              reg647 = $unsigned((reg583 ?
                  ($unsigned((~|reg494)) || {(reg518 ?
                          (8'ha2) : reg602)}) : (~|(&$unsigned(reg592)))));
              reg651 = {($unsigned($unsigned(reg595[(4'hf):(3'h7)])) ?
                      $unsigned(reg501) : ($signed((^reg626)) ?
                          ((~reg645) <= (-reg551)) : reg623)),
                  reg481};
              reg653 <= $unsigned($signed($signed(reg553)));
            end
        end
      reg654 = reg501;
      reg655 = (~((|reg606[(2'h3):(1'h1)]) ?
          reg521[(4'ha):(4'ha)] : $signed($signed(((8'h9f) ~^ reg510)))));
    end
  always
    @(posedge clk) begin
      for (forvar656 = (1'h0); (forvar656 < (2'h3)); forvar656 = (forvar656 + (1'h1)))
        begin
          reg657 <= reg600[(2'h3):(1'h1)];
          reg658 <= ((7'h41) > reg494);
          for (forvar659 = (1'h0); (forvar659 < (1'h0)); forvar659 = (forvar659 + (1'h1)))
            begin
              reg660 <= ($signed({$signed($signed((8'hb2)))}) ?
                  (~reg544) : reg544);
              reg661 = (&reg613[(4'h8):(4'h8)]);
              reg662 <= reg648;
            end
          if (($unsigned((reg613 ?
              reg560[(3'h4):(2'h2)] : reg642[(1'h0):(1'h0)])) ^~ (!(8'hab))))
            begin
              reg663 = $unsigned($signed(reg571[(4'hb):(2'h2)]));
              reg664 = (reg476[(1'h0):(1'h0)] | $signed(reg627[(1'h1):(1'h1)]));
              reg665 <= (($unsigned($signed($unsigned(reg658))) ?
                  $signed($unsigned($unsigned(reg661))) : (reg543 && (reg629 ?
                      (8'h9e) : (reg500 ^ wire471)))) | (reg561[(3'h6):(3'h6)] >>> ($unsigned($unsigned(reg488)) ~^ (reg611 ?
                  reg623 : (^~reg517)))));
            end
          else
            begin
              reg665 <= (+{(|(reg478 ? (reg648 | reg569) : $unsigned((8'h9e)))),
                  reg605});
              reg666 <= ((^~($unsigned($unsigned(reg615)) << ({reg643,
                      reg488} & reg569))) ?
                  $unsigned((~reg508)) : reg474[(4'he):(2'h2)]);
              reg667 <= ((8'hbf) > (!reg585));
              reg668 <= (reg661 <<< reg627);
            end
        end
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module72  (y, clk, wire73, wire74, wire75, wire76);
  output wire [(32'h28f):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire73;
  input wire signed [(5'h12):(1'h0)] wire74;
  input wire [(5'h10):(1'h0)] wire75;
  input wire signed [(4'hc):(1'h0)] wire76;
  wire signed [(5'h14):(1'h0)] wire431;
  wire signed [(3'h7):(1'h0)] wire275;
  wire [(5'h11):(1'h0)] wire95;
  wire signed [(4'hc):(1'h0)] wire273;
  reg [(5'h11):(1'h0)] reg459 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg458 = (1'h0);
  reg [(4'hf):(1'h0)] reg457 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg456 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg454 = (1'h0);
  reg [(4'hb):(1'h0)] reg453 = (1'h0);
  reg [(4'hf):(1'h0)] reg450 = (1'h0);
  reg [(3'h7):(1'h0)] reg448 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg446 = (1'h0);
  reg [(5'h10):(1'h0)] reg445 = (1'h0);
  reg [(5'h11):(1'h0)] reg444 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg443 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg442 = (1'h0);
  reg [(2'h3):(1'h0)] reg440 = (1'h0);
  reg [(5'h12):(1'h0)] reg438 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg437 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg436 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg435 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg434 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg80 = (1'h0);
  reg [(5'h10):(1'h0)] reg81 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg86 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg89 = (1'h0);
  reg [(4'hb):(1'h0)] reg90 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg93 = (1'h0);
  reg [(3'h4):(1'h0)] reg94 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg460 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg455 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg452 = (1'h0);
  reg [(2'h2):(1'h0)] reg451 = (1'h0);
  reg [(5'h10):(1'h0)] forvar449 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar447 = (1'h0);
  reg [(5'h15):(1'h0)] reg441 = (1'h0);
  reg [(5'h12):(1'h0)] forvar434 = (1'h0);
  reg [(4'ha):(1'h0)] reg439 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg433 = (1'h0);
  reg signed [(4'he):(1'h0)] reg92 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg91 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg88 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg87 = (1'h0);
  reg signed [(4'he):(1'h0)] reg85 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar84 = (1'h0);
  reg [(4'hf):(1'h0)] reg83 = (1'h0);
  reg [(5'h11):(1'h0)] reg82 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg79 = (1'h0);
  reg [(4'he):(1'h0)] forvar78 = (1'h0);
  reg [(3'h4):(1'h0)] forvar77 = (1'h0);
  assign y = {wire431,
                 wire275,
                 wire95,
                 wire273,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg454,
                 reg453,
                 reg450,
                 reg448,
                 reg446,
                 reg445,
                 reg444,
                 reg443,
                 reg442,
                 reg440,
                 reg438,
                 reg437,
                 reg436,
                 reg435,
                 reg434,
                 reg80,
                 reg81,
                 reg86,
                 reg89,
                 reg90,
                 reg93,
                 reg94,
                 reg460,
                 reg455,
                 reg452,
                 reg451,
                 forvar449,
                 forvar447,
                 reg441,
                 forvar434,
                 reg439,
                 reg433,
                 reg92,
                 reg91,
                 reg88,
                 reg87,
                 reg85,
                 forvar84,
                 reg83,
                 reg82,
                 reg79,
                 forvar78,
                 forvar77,
                 (1'h0)};
  always
    @(posedge clk) begin
      for (forvar77 = (1'h0); (forvar77 < (1'h0)); forvar77 = (forvar77 + (1'h1)))
        begin
          for (forvar78 = (1'h0); (forvar78 < (1'h1)); forvar78 = (forvar78 + (1'h1)))
            begin
              reg79 = {($unsigned((8'hb6)) ? (8'hb7) : (~wire76)),
                  ($signed((wire73[(4'h9):(2'h2)] ?
                          wire75[(4'ha):(3'h4)] : ((8'hba) ?
                              wire74 : forvar77))) ?
                      (((forvar77 ? wire76 : wire74) == wire73[(4'hd):(3'h6)]) ?
                          (^~(wire73 << (7'h42))) : $signed(wire73)) : (wire74[(4'he):(3'h4)] >= wire74[(1'h0):(1'h0)]))};
              reg80 <= (~((^({forvar77} == $unsigned((8'had)))) || $signed($signed((wire76 ?
                  wire76 : forvar78)))));
              reg81 <= (wire76 ?
                  (forvar78[(2'h3):(2'h2)] ?
                      (wire76[(3'h6):(3'h6)] != forvar78) : reg80[(2'h3):(2'h3)]) : $unsigned(forvar77[(2'h3):(1'h0)]));
            end
          reg82 = wire73[(5'h12):(3'h6)];
        end
      reg83 = ({wire75} < $unsigned(((reg82[(2'h2):(1'h0)] ?
          (~(7'h42)) : reg80[(2'h3):(1'h0)]) * reg79)));
      for (forvar84 = (1'h0); (forvar84 < (1'h0)); forvar84 = (forvar84 + (1'h1)))
        begin
          reg85 = reg83[(4'he):(3'h4)];
          reg86 <= (wire73 ?
              (($unsigned($signed((8'ha6))) ? reg79 : {$signed(reg83)}) ?
                  $unsigned($signed(reg83)) : (forvar78[(4'hc):(4'hb)] ?
                      (~^(reg80 ?
                          reg81 : (8'ha0))) : reg83[(4'hf):(3'h7)])) : reg80);
          if ((reg82 ?
              $signed(($unsigned((wire73 <<< reg81)) ?
                  reg81[(4'h8):(4'h8)] : forvar78[(4'he):(3'h6)])) : wire75))
            begin
              reg87 = forvar84;
              reg88 = {reg83};
              reg89 <= wire75[(4'hb):(4'ha)];
              reg90 <= wire73;
            end
          else
            begin
              reg89 <= wire76;
              reg91 = $unsigned(wire73);
              reg92 = forvar84;
            end
          reg93 <= ({reg91} && ((8'ha1) ?
              (+reg92[(2'h2):(1'h1)]) : {wire75[(4'hd):(4'ha)]}));
        end
      reg94 <= reg79[(3'h6):(3'h5)];
    end
  assign wire95 = ((^{reg86, $signed($unsigned(reg94))}) ?
                      (wire73[(3'h7):(2'h2)] ?
                          {$unsigned((wire76 * (8'hab))),
                              {$signed(reg89)}} : $signed({(^wire75),
                              reg81[(4'h8):(4'h8)]})) : $unsigned((^~(((8'hae) >= reg90) ?
                          {reg80, (8'h9f)} : wire73))));
  module96 #() modinst274 (.wire99(wire74), .wire101(wire95), .wire97(wire73), .y(wire273), .wire100(reg89), .wire98(reg86), .clk(clk));
  assign wire275 = ({$signed((!(wire74 - wire273)))} - wire73[(3'h6):(1'h0)]);
  module276 #() modinst432 (wire431, clk, reg80, wire73, wire75, reg94, reg90);
  always
    @(posedge clk) begin
      if (((8'hac) ?
          $signed($signed((-wire273))) : $unsigned(((|wire275) ?
              wire75[(4'ha):(4'h8)] : (+reg81)))))
        begin
          if (($signed($signed(reg93[(5'h10):(4'hf)])) ?
              $signed(((wire431[(3'h6):(2'h2)] ?
                  ((8'hbb) ?
                      wire95 : reg81) : (+reg81)) != wire431[(3'h4):(2'h3)])) : reg89[(1'h0):(1'h0)]))
            begin
              reg433 = wire95;
              reg434 <= $unsigned((-($signed(wire76) ?
                  $signed((8'hb0)) : (-$signed(reg80)))));
              reg435 <= wire73;
              reg436 <= $unsigned((+($unsigned(wire273) ?
                  ((wire76 ? wire95 : wire275) ?
                      $unsigned(reg435) : $signed(wire273)) : (8'hae))));
              reg437 <= (reg433[(1'h0):(1'h0)] ?
                  {(wire95 ? wire275 : reg80[(3'h7):(2'h3)]),
                      $unsigned(({reg94, reg80} ?
                          wire273[(1'h1):(1'h1)] : $unsigned((8'hb2))))} : wire74[(1'h0):(1'h0)]);
            end
          else
            begin
              reg434 <= (reg437 ?
                  {(reg437 & $signed($signed((8'hbe)))),
                      reg93} : $unsigned($signed(reg80)));
              reg435 <= $unsigned(wire73);
              reg436 <= (7'h41);
              reg437 <= $unsigned($signed((~^(~|(&reg80)))));
              reg438 <= reg435[(3'h4):(1'h1)];
            end
          reg439 = $signed(reg94);
        end
      else
        begin
          reg433 = (&$unsigned(($unsigned({wire74, reg436}) ?
              reg80 : wire431[(3'h4):(3'h4)])));
          for (forvar434 = (1'h0); (forvar434 < (2'h2)); forvar434 = (forvar434 + (1'h1)))
            begin
              reg439 = (-$unsigned(reg439));
            end
          if ((~&$unsigned($unsigned((!{reg433})))))
            begin
              reg440 <= (~((-({reg80} ^ $unsigned(reg89))) && $signed((~&reg93[(1'h1):(1'h1)]))));
              reg441 = $signed(reg435);
            end
          else
            begin
              reg440 <= (reg441 ?
                  ((^~(wire74 >>> $unsigned(forvar434))) ?
                      reg435[(3'h5):(1'h1)] : reg434[(4'h8):(4'h8)]) : $signed((({reg86,
                          wire95} ?
                      forvar434 : (wire431 ?
                          wire95 : wire73)) >>> (reg439 < (8'hae)))));
              reg442 <= reg438;
              reg443 <= $unsigned(wire431);
              reg444 <= (~($signed((wire74[(1'h0):(1'h0)] + reg80)) >= wire75));
              reg445 <= wire431;
            end
          reg446 <= reg86[(4'ha):(3'h4)];
        end
      for (forvar447 = (1'h0); (forvar447 < (1'h0)); forvar447 = (forvar447 + (1'h1)))
        begin
          reg448 <= $unsigned($signed(($unsigned(reg86[(1'h1):(1'h0)]) | (((8'hba) ^~ wire273) ?
              $unsigned(wire95) : (+reg86)))));
          for (forvar449 = (1'h0); (forvar449 < (1'h1)); forvar449 = (forvar449 + (1'h1)))
            begin
              reg450 <= (^(!(~^$signed(reg94))));
              reg451 = reg448[(3'h7):(3'h4)];
              reg452 = $unsigned((reg433 ?
                  ($unsigned($signed((8'ha9))) ?
                      wire75 : forvar447[(2'h3):(2'h2)]) : $signed((reg80[(1'h1):(1'h0)] ?
                      (~|forvar449) : {forvar449, wire75}))));
              reg453 <= (reg442[(3'h6):(2'h2)] ? reg90 : $unsigned(wire275));
            end
        end
    end
  always
    @(posedge clk) begin
      reg454 <= reg448[(3'h7):(1'h1)];
      reg455 = reg90;
      reg456 <= reg81[(4'he):(4'hc)];
      reg457 <= reg455[(3'h6):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg458 <= (8'ha6);
      reg459 <= $signed($unsigned($unsigned($unsigned((^~reg458)))));
      reg460 = (reg86 || (reg438 ? wire431 : $unsigned((~&$unsigned(reg440)))));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module276
#(parameter param429 = ((8'hb2) ? (8'hbc) : ((-{((8'hbf) & (8'ha7)), ((7'h41) ^ (8'hac))}) || {(((8'hb4) || (8'ha7)) == ((8'h9d) != (8'ha6))), (((7'h41) ? (8'haf) : (8'ha1)) ? ((8'h9f) != (8'ha8)) : ((8'hb8) ? (8'hb8) : (8'h9f)))})), 
parameter param430 = (~&(((~param429) ? param429 : ((param429 ? param429 : param429) > (&param429))) ? (((^~(8'hbe)) ? (~^param429) : (param429 ? param429 : param429)) > param429) : ((~|(param429 <<< param429)) & (param429 ~^ param429)))))
(y, clk, wire281, wire280, wire279, wire278, wire277);
  output wire [(32'h72a):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h11):(1'h0)] wire281;
  input wire signed [(4'hf):(1'h0)] wire280;
  input wire signed [(5'h10):(1'h0)] wire279;
  input wire [(3'h4):(1'h0)] wire278;
  input wire [(4'hb):(1'h0)] wire277;
  wire signed [(3'h7):(1'h0)] wire420;
  wire signed [(4'hf):(1'h0)] wire319;
  reg signed [(3'h6):(1'h0)] reg428 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg427 = (1'h0);
  reg [(4'hc):(1'h0)] reg425 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg422 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg419 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg418 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg416 = (1'h0);
  reg [(4'hf):(1'h0)] reg414 = (1'h0);
  reg [(5'h15):(1'h0)] reg412 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg411 = (1'h0);
  reg [(5'h12):(1'h0)] reg410 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg409 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg407 = (1'h0);
  reg [(4'ha):(1'h0)] reg406 = (1'h0);
  reg signed [(4'he):(1'h0)] reg405 = (1'h0);
  reg [(2'h2):(1'h0)] reg402 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg401 = (1'h0);
  reg [(3'h6):(1'h0)] reg398 = (1'h0);
  reg [(3'h6):(1'h0)] reg396 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg394 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg393 = (1'h0);
  reg [(3'h6):(1'h0)] reg392 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg389 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg388 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg387 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg385 = (1'h0);
  reg [(4'he):(1'h0)] reg381 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg379 = (1'h0);
  reg signed [(4'he):(1'h0)] reg378 = (1'h0);
  reg [(5'h15):(1'h0)] reg376 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg375 = (1'h0);
  reg [(5'h11):(1'h0)] reg374 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg373 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg372 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg371 = (1'h0);
  reg [(5'h10):(1'h0)] reg369 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg367 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg365 = (1'h0);
  reg [(5'h14):(1'h0)] reg359 = (1'h0);
  reg [(2'h3):(1'h0)] reg358 = (1'h0);
  reg [(4'hd):(1'h0)] reg357 = (1'h0);
  reg [(3'h6):(1'h0)] reg355 = (1'h0);
  reg [(5'h10):(1'h0)] reg354 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg351 = (1'h0);
  reg [(3'h4):(1'h0)] reg348 = (1'h0);
  reg [(5'h14):(1'h0)] reg345 = (1'h0);
  reg [(4'hb):(1'h0)] reg341 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg342 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg336 = (1'h0);
  reg [(2'h2):(1'h0)] reg330 = (1'h0);
  reg [(2'h2):(1'h0)] reg340 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg339 = (1'h0);
  reg [(2'h3):(1'h0)] reg337 = (1'h0);
  reg [(4'h9):(1'h0)] reg334 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg332 = (1'h0);
  reg [(4'h9):(1'h0)] reg331 = (1'h0);
  reg [(2'h3):(1'h0)] reg327 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg326 = (1'h0);
  reg [(5'h11):(1'h0)] reg324 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg321 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg320 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg317 = (1'h0);
  reg [(5'h15):(1'h0)] reg315 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg314 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg309 = (1'h0);
  reg [(4'hd):(1'h0)] reg308 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg306 = (1'h0);
  reg [(5'h10):(1'h0)] reg305 = (1'h0);
  reg [(5'h11):(1'h0)] reg304 = (1'h0);
  reg [(4'hf):(1'h0)] reg303 = (1'h0);
  reg [(3'h5):(1'h0)] reg301 = (1'h0);
  reg [(5'h11):(1'h0)] reg299 = (1'h0);
  reg [(4'ha):(1'h0)] reg297 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg296 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg295 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg292 = (1'h0);
  reg signed [(4'he):(1'h0)] reg289 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg288 = (1'h0);
  reg [(4'ha):(1'h0)] reg287 = (1'h0);
  reg [(4'h8):(1'h0)] reg286 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg285 = (1'h0);
  reg [(4'he):(1'h0)] reg284 = (1'h0);
  reg [(3'h4):(1'h0)] reg426 = (1'h0);
  reg [(4'hb):(1'h0)] reg424 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar423 = (1'h0);
  reg [(5'h10):(1'h0)] forvar421 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg417 = (1'h0);
  reg [(2'h3):(1'h0)] forvar415 = (1'h0);
  reg [(3'h5):(1'h0)] forvar413 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar408 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg404 = (1'h0);
  reg [(4'h9):(1'h0)] reg403 = (1'h0);
  reg [(4'hd):(1'h0)] forvar400 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg399 = (1'h0);
  reg [(4'hd):(1'h0)] reg397 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar395 = (1'h0);
  reg [(4'hc):(1'h0)] reg391 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg390 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg386 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg384 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar383 = (1'h0);
  reg [(3'h6):(1'h0)] forvar382 = (1'h0);
  reg [(3'h7):(1'h0)] reg380 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar377 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar370 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg368 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg366 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg364 = (1'h0);
  reg [(4'hc):(1'h0)] reg363 = (1'h0);
  reg [(5'h14):(1'h0)] reg362 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar361 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg360 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar356 = (1'h0);
  reg [(3'h6):(1'h0)] forvar353 = (1'h0);
  reg [(3'h5):(1'h0)] forvar352 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg350 = (1'h0);
  reg [(2'h3):(1'h0)] reg349 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg347 = (1'h0);
  reg [(5'h11):(1'h0)] forvar346 = (1'h0);
  reg [(4'hf):(1'h0)] forvar342 = (1'h0);
  reg [(5'h13):(1'h0)] reg344 = (1'h0);
  reg [(4'hc):(1'h0)] reg343 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar341 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar331 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg338 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar336 = (1'h0);
  reg [(4'hf):(1'h0)] reg335 = (1'h0);
  reg [(5'h12):(1'h0)] reg333 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar330 = (1'h0);
  reg [(4'h8):(1'h0)] reg329 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg328 = (1'h0);
  reg [(5'h13):(1'h0)] reg325 = (1'h0);
  reg [(2'h3):(1'h0)] reg323 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg322 = (1'h0);
  reg [(5'h14):(1'h0)] reg318 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg316 = (1'h0);
  reg [(3'h4):(1'h0)] reg313 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar311 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg310 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg307 = (1'h0);
  reg [(3'h6):(1'h0)] reg302 = (1'h0);
  reg [(3'h7):(1'h0)] forvar300 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar298 = (1'h0);
  reg [(4'hb):(1'h0)] reg294 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg293 = (1'h0);
  reg [(3'h5):(1'h0)] reg291 = (1'h0);
  reg [(4'hc):(1'h0)] forvar291 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg290 = (1'h0);
  reg [(4'hb):(1'h0)] forvar283 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg282 = (1'h0);
  assign y = {wire420,
                 wire319,
                 reg428,
                 reg427,
                 reg425,
                 reg422,
                 reg419,
                 reg418,
                 reg416,
                 reg414,
                 reg412,
                 reg411,
                 reg410,
                 reg409,
                 reg407,
                 reg406,
                 reg405,
                 reg402,
                 reg401,
                 reg398,
                 reg396,
                 reg394,
                 reg393,
                 reg392,
                 reg389,
                 reg388,
                 reg387,
                 reg385,
                 reg381,
                 reg379,
                 reg378,
                 reg376,
                 reg375,
                 reg374,
                 reg373,
                 reg372,
                 reg371,
                 reg369,
                 reg367,
                 reg365,
                 reg359,
                 reg358,
                 reg357,
                 reg355,
                 reg354,
                 reg351,
                 reg348,
                 reg345,
                 reg341,
                 reg342,
                 reg336,
                 reg330,
                 reg340,
                 reg339,
                 reg337,
                 reg334,
                 reg332,
                 reg331,
                 reg327,
                 reg326,
                 reg324,
                 reg321,
                 reg320,
                 reg317,
                 reg315,
                 reg314,
                 reg312,
                 reg309,
                 reg308,
                 reg306,
                 reg305,
                 reg304,
                 reg303,
                 reg301,
                 reg299,
                 reg297,
                 reg296,
                 reg295,
                 reg292,
                 reg289,
                 reg288,
                 reg287,
                 reg286,
                 reg285,
                 reg284,
                 reg426,
                 reg424,
                 forvar423,
                 forvar421,
                 reg417,
                 forvar415,
                 forvar413,
                 forvar408,
                 reg404,
                 reg403,
                 forvar400,
                 reg399,
                 reg397,
                 forvar395,
                 reg391,
                 reg390,
                 reg386,
                 reg384,
                 forvar383,
                 forvar382,
                 reg380,
                 forvar377,
                 forvar370,
                 reg368,
                 reg366,
                 reg364,
                 reg363,
                 reg362,
                 forvar361,
                 reg360,
                 forvar356,
                 forvar353,
                 forvar352,
                 reg350,
                 reg349,
                 reg347,
                 forvar346,
                 forvar342,
                 reg344,
                 reg343,
                 forvar341,
                 forvar331,
                 reg338,
                 forvar336,
                 reg335,
                 reg333,
                 forvar330,
                 reg329,
                 reg328,
                 reg325,
                 reg323,
                 reg322,
                 reg318,
                 reg316,
                 reg313,
                 forvar311,
                 reg310,
                 reg307,
                 reg302,
                 forvar300,
                 forvar298,
                 reg294,
                 reg293,
                 reg291,
                 forvar291,
                 reg290,
                 forvar283,
                 reg282,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg282 = (7'h44);
    end
  always
    @(posedge clk) begin
      for (forvar283 = (1'h0); (forvar283 < (3'h4)); forvar283 = (forvar283 + (1'h1)))
        begin
          if ($unsigned($unsigned($signed(wire280))))
            begin
              reg284 <= (wire279 ?
                  ({{(wire279 ?
                              (8'h9d) : (7'h42))}} >>> wire277[(2'h3):(2'h3)]) : (wire279[(4'hf):(3'h4)] ?
                      (wire281[(4'h9):(3'h4)] & $unsigned((wire277 | wire277))) : {((~&wire278) ?
                              $signed(wire281) : wire281[(4'h8):(1'h0)])}));
              reg285 <= wire278[(2'h3):(2'h2)];
            end
          else
            begin
              reg284 <= (($unsigned(((forvar283 ?
                  wire280 : wire278) >> $signed(wire279))) ~^ wire279) | {$signed($signed(wire277[(3'h4):(2'h3)])),
                  $unsigned(reg284[(4'he):(4'ha)])});
              reg285 <= $unsigned($signed((reg285 >>> wire277)));
            end
          reg286 <= (wire279 ^ $signed((~&(^(^wire280)))));
          reg287 <= reg286;
          reg288 <= {(reg285[(1'h1):(1'h0)] ?
                  (-$unsigned((-wire281))) : $signed(($unsigned(wire280) * $signed((8'hb8)))))};
        end
      if ((({wire277[(1'h1):(1'h1)]} ?
          $signed((~wire278)) : reg287[(4'h9):(1'h0)]) * {{reg287[(1'h1):(1'h0)]}}))
        begin
          reg289 <= $signed(($signed((-$signed(forvar283))) <= $signed($signed(reg288[(3'h4):(3'h4)]))));
          reg290 = $unsigned(reg285[(4'h9):(3'h7)]);
          for (forvar291 = (1'h0); (forvar291 < (3'h4)); forvar291 = (forvar291 + (1'h1)))
            begin
              reg292 <= {(&wire277[(3'h6):(3'h4)]),
                  $unsigned(({reg284, reg286} ^ ((forvar283 ?
                      forvar283 : (8'ha3)) != {reg288})))};
            end
        end
      else
        begin
          if ((($unsigned((wire278[(1'h0):(1'h0)] ?
                  ((8'ha3) ?
                      reg290 : (8'hba)) : $unsigned(reg290))) + {reg292[(4'hb):(3'h4)],
                  $unsigned((!wire280))}) ?
              ((&((reg292 ?
                  wire281 : forvar291) << wire280)) >>> forvar291[(3'h4):(3'h4)]) : $signed((-reg287[(1'h0):(1'h0)]))))
            begin
              reg290 = reg292[(2'h3):(2'h2)];
              reg291 = (((reg287[(2'h3):(1'h1)] ~^ ($unsigned(forvar283) ?
                      $unsigned((8'hac)) : (wire277 >> reg286))) - wire279[(4'hc):(1'h1)]) ?
                  ((((~reg286) && wire279) ? (8'ha7) : reg288[(1'h0):(1'h0)]) ?
                      $signed(((+reg289) ^~ reg289)) : reg287[(1'h0):(1'h0)]) : {(&$signed($unsigned(reg285)))});
              reg293 = {(~^$unsigned((8'hae)))};
              reg294 = $unsigned(((&(|$unsigned(reg285))) ?
                  (~|reg286) : reg288));
              reg295 <= forvar291[(3'h5):(2'h3)];
            end
          else
            begin
              reg289 <= (wire277[(3'h7):(1'h1)] ?
                  $signed(reg295) : $unsigned($unsigned((~^{reg290,
                      forvar283}))));
              reg292 <= reg284[(3'h7):(3'h6)];
            end
          reg296 <= $signed(reg288);
          reg297 <= $signed((~|{($unsigned(wire278) >> (^reg296)),
              reg296[(2'h3):(1'h0)]}));
        end
      for (forvar298 = (1'h0); (forvar298 < (2'h2)); forvar298 = (forvar298 + (1'h1)))
        begin
          reg299 <= $signed(reg290[(3'h5):(2'h2)]);
          for (forvar300 = (1'h0); (forvar300 < (2'h2)); forvar300 = (forvar300 + (1'h1)))
            begin
              reg301 <= reg288[(3'h6):(3'h4)];
              reg302 = $unsigned({reg296[(3'h6):(1'h1)]});
              reg303 <= ((~^(reg292[(4'hc):(3'h4)] ?
                  (8'hb9) : forvar300[(1'h1):(1'h1)])) == forvar300);
            end
          if ($unsigned((({(8'hb8)} ?
              ({reg294,
                  reg303} ~^ forvar291) : reg287[(1'h1):(1'h0)]) ^~ (~|{(wire278 && forvar291),
              (-wire281)}))))
            begin
              reg304 <= (reg303 ? wire279 : {$signed((^reg293)), forvar298});
              reg305 <= $signed($unsigned((reg293[(1'h0):(1'h0)] >>> {reg292[(1'h0):(1'h0)],
                  (8'hbe)})));
              reg306 <= {(-$signed(wire279[(4'h8):(3'h7)])),
                  (|{$signed((wire280 ? forvar300 : reg287)),
                      (reg304 <<< {reg296})})};
            end
          else
            begin
              reg304 <= ($signed((~^reg291)) ? reg293[(2'h2):(1'h0)] : reg285);
              reg307 = ((^~$unsigned(($signed(reg299) <= ((8'h9d) ?
                  wire277 : forvar291)))) ^ (~&$unsigned($signed((reg297 * (8'h9c))))));
              reg308 <= $signed((((wire281 ?
                  reg304 : reg284[(2'h2):(1'h1)]) <<< $signed(reg292[(4'ha):(4'ha)])) * (reg306[(3'h5):(3'h5)] ?
                  reg296 : (~&(reg303 + (8'hb0))))));
              reg309 <= (reg305[(4'he):(4'h8)] >> {$signed($unsigned((8'hb2)))});
              reg310 = $signed(reg289[(4'h9):(2'h3)]);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar311 = (1'h0); (forvar311 < (3'h4)); forvar311 = (forvar311 + (1'h1)))
        begin
          reg312 <= reg306[(2'h2):(1'h0)];
        end
      reg313 = (reg286 * reg296[(1'h0):(1'h0)]);
      reg314 <= ((~^forvar311) ? reg285 : (~|reg303[(3'h6):(3'h6)]));
      reg315 <= $unsigned((^~$signed(reg292[(1'h0):(1'h0)])));
    end
  always
    @(posedge clk) begin
      reg316 = (&$signed(reg304));
      reg317 <= reg314;
      reg318 = reg306;
    end
  assign wire319 = ((~|(^~(-$signed(reg306)))) ?
                       $unsigned((&wire281)) : {$unsigned(reg286[(3'h5):(1'h0)])});
  always
    @(posedge clk) begin
      reg320 <= ((((+((8'hb5) ? reg284 : (8'ha1))) ?
              ((reg295 ?
                  reg309 : (8'had)) != ((8'hbe) | reg288)) : (reg295[(3'h5):(2'h3)] ?
                  {reg299, (7'h41)} : ((8'ha0) ?
                      reg289 : reg304))) | ($unsigned(wire277[(3'h7):(3'h7)]) ^~ (~{reg297,
              reg315}))) ?
          reg303 : ({reg286[(1'h1):(1'h0)]} ?
              {wire319[(2'h3):(1'h0)],
                  ($signed((8'hac)) ?
                      reg303 : {reg301, reg292})} : reg295[(3'h4):(1'h0)]));
      reg321 <= (~|reg312[(1'h0):(1'h0)]);
    end
  always
    @(posedge clk) begin
      reg322 = ($unsigned((^~(~$signed((8'ha4))))) ?
          (^~({reg304, reg284} + {reg312[(4'hd):(4'ha)],
              (reg287 ? reg296 : reg286)})) : (~|{reg299[(1'h0):(1'h0)],
              wire281}));
    end
  always
    @(posedge clk) begin
      reg323 = reg289[(3'h5):(1'h0)];
      reg324 <= $signed((~&wire319[(3'h7):(1'h1)]));
      reg325 = (reg320 && reg309);
      reg326 <= reg284;
    end
  always
    @(posedge clk) begin
      reg327 <= $unsigned($signed($unsigned({(wire277 < reg312),
          reg314[(1'h1):(1'h0)]})));
    end
  always
    @(posedge clk) begin
      if ($unsigned(($signed($signed((wire277 ?
          reg287 : reg289))) && (~^$signed((reg315 & reg315))))))
        begin
          reg328 = reg301[(1'h0):(1'h0)];
          reg329 = (+$unsigned((~&reg304[(5'h10):(4'he)])));
          for (forvar330 = (1'h0); (forvar330 < (2'h2)); forvar330 = (forvar330 + (1'h1)))
            begin
              reg331 <= reg287[(3'h6):(3'h4)];
              reg332 <= ({{({reg292} ^ reg301)}} >= {($signed((reg305 ?
                          wire277 : reg328)) ?
                      $unsigned($signed(wire280)) : ($signed(reg320) ^~ reg297[(2'h3):(2'h3)]))});
              reg333 = {($signed(reg288[(1'h0):(1'h0)]) ?
                      wire277 : reg305[(1'h1):(1'h1)])};
              reg334 <= ($signed(($unsigned(reg305) ?
                      reg292 : ($signed(reg284) ?
                          (reg299 | (8'hae)) : reg285[(3'h7):(3'h5)]))) ?
                  (reg306 ?
                      (((~|reg320) >>> $signed(reg288)) ?
                          (~$unsigned(reg309)) : reg286) : wire280) : $signed($signed(wire280[(4'h9):(1'h1)])));
              reg335 = (+{wire281[(3'h6):(2'h3)]});
            end
          for (forvar336 = (1'h0); (forvar336 < (2'h2)); forvar336 = (forvar336 + (1'h1)))
            begin
              reg337 <= {reg296};
              reg338 = reg288[(1'h0):(1'h0)];
              reg339 <= (|$unsigned(($signed(((8'hbd) ? reg292 : reg306)) ?
                  ($unsigned((8'ha5)) < (wire279 ?
                      (8'hb1) : reg335)) : $signed($signed(reg333)))));
              reg340 <= $signed(({reg284[(3'h7):(2'h3)],
                  ($signed(reg337) ?
                      (reg315 << reg287) : reg332)} ~^ {wire281[(4'ha):(4'h9)],
                  (+(reg284 ? reg312 : reg328))}));
            end
        end
      else
        begin
          reg330 <= $signed(reg337[(2'h2):(1'h1)]);
          for (forvar331 = (1'h0); (forvar331 < (2'h2)); forvar331 = (forvar331 + (1'h1)))
            begin
              reg333 = (~({{(~|reg289)}, (reg304 | $signed(reg299))} ?
                  reg334 : ((((8'hbf) << reg308) - $unsigned(reg314)) <= (reg285 & $signed(reg321)))));
              reg335 = (({$unsigned((reg315 ? (8'hab) : reg308)),
                          ($signed((8'hb2)) ? (~&reg304) : $unsigned(reg314))} ?
                      $unsigned(reg324[(2'h3):(2'h3)]) : $unsigned((+(reg309 >>> reg308)))) ?
                  $signed({((reg286 ? reg320 : forvar336) ?
                          {reg337} : ((8'hbc) ?
                              wire279 : wire278))}) : {$signed((+wire280))});
              reg336 <= $signed(reg299[(5'h10):(4'h8)]);
            end
        end
      if ($signed((forvar336[(4'h9):(4'h9)] ?
          reg331[(1'h1):(1'h0)] : $unsigned({(reg320 ? forvar336 : reg285),
              (reg337 >> reg336)}))))
        begin
          for (forvar341 = (1'h0); (forvar341 < (3'h4)); forvar341 = (forvar341 + (1'h1)))
            begin
              reg342 <= reg309;
              reg343 = reg292[(5'h11):(4'h8)];
            end
          reg344 = forvar341[(2'h3):(2'h2)];
        end
      else
        begin
          reg341 <= (forvar336[(3'h4):(1'h1)] ?
              ((~^$unsigned((reg336 <<< reg317))) ?
                  $unsigned(($unsigned(reg288) ?
                      reg315[(4'hd):(4'hb)] : (reg337 ?
                          reg306 : reg334))) : reg314[(1'h0):(1'h0)]) : ($signed(wire281[(4'hf):(3'h4)]) < $signed((^(reg304 - wire279)))));
          for (forvar342 = (1'h0); (forvar342 < (1'h0)); forvar342 = (forvar342 + (1'h1)))
            begin
              reg345 <= reg328;
            end
        end
      for (forvar346 = (1'h0); (forvar346 < (2'h2)); forvar346 = (forvar346 + (1'h1)))
        begin
          reg347 = reg321[(2'h3):(1'h0)];
          reg348 <= ((~^reg306) | (($signed(reg285[(2'h2):(2'h2)]) ?
              $unsigned((&reg329)) : (8'ha1)) >= $signed((8'ha5))));
          reg349 = reg320;
          reg350 = $signed($signed({($unsigned(wire278) ?
                  $signed((8'ha3)) : {reg301, (7'h41)}),
              (&$unsigned(reg303))}));
          reg351 <= ($signed((reg344 == $unsigned(reg329))) ~^ reg320[(3'h5):(3'h5)]);
        end
      for (forvar352 = (1'h0); (forvar352 < (1'h0)); forvar352 = (forvar352 + (1'h1)))
        begin
          for (forvar353 = (1'h0); (forvar353 < (2'h2)); forvar353 = (forvar353 + (1'h1)))
            begin
              reg354 <= $signed((+$signed(reg337[(1'h1):(1'h0)])));
            end
          reg355 <= $signed((-({(7'h44), forvar331[(4'hd):(1'h0)]} ?
              reg297 : (~|(reg284 ? (8'haf) : reg296)))));
          for (forvar356 = (1'h0); (forvar356 < (1'h0)); forvar356 = (forvar356 + (1'h1)))
            begin
              reg357 <= ((((+(reg341 - reg306)) && (reg344 ?
                      $signed(reg292) : $signed(reg308))) ?
                  reg344 : $signed($unsigned((reg342 ?
                      reg339 : (7'h41))))) >> (reg312[(4'h9):(3'h4)] ?
                  (~&wire279[(4'h8):(3'h7)]) : reg327));
            end
          reg358 <= forvar336[(4'ha):(4'h8)];
          reg359 <= (wire279[(4'hb):(2'h3)] ?
              wire278 : {$signed({{reg337, reg340}, (~&(8'h9d))})});
        end
    end
  always
    @(posedge clk) begin
      reg360 = ($unsigned(({(reg330 ~^ wire281)} ?
              ($signed(reg305) ?
                  (reg303 ?
                      reg317 : reg309) : $signed(reg297)) : (reg345[(3'h7):(3'h5)] ?
                  $unsigned(reg314) : $unsigned(reg306)))) ?
          {($unsigned(reg334) ?
                  $unsigned((reg354 ?
                      reg348 : (8'ha1))) : ((7'h44) << (!reg359)))} : reg351);
      for (forvar361 = (1'h0); (forvar361 < (1'h1)); forvar361 = (forvar361 + (1'h1)))
        begin
          reg362 = ((~($unsigned((8'hb4)) ?
                  reg305[(1'h1):(1'h0)] : (reg351 ?
                      $unsigned(reg284) : $unsigned(wire277)))) ?
              (+({reg327} < $signed(reg309))) : reg285[(3'h7):(2'h3)]);
        end
      reg363 = $signed({{$unsigned($unsigned((8'ha5))),
              ($unsigned(reg336) ? (~reg301) : $unsigned(reg303))},
          $unsigned(reg317)});
      reg364 = reg320[(4'hf):(4'h9)];
    end
  always
    @(posedge clk) begin
      if (reg330[(2'h2):(1'h0)])
        begin
          reg365 <= $unsigned(reg357[(4'h9):(2'h2)]);
        end
      else
        begin
          reg366 = (+(reg309 ?
              reg331 : ($unsigned((wire280 ? reg337 : wire279)) + reg337)));
          reg367 <= reg295;
          reg368 = reg297[(3'h5):(3'h4)];
          reg369 <= (reg314[(1'h1):(1'h1)] ?
              (reg341 ?
                  $signed(reg339[(3'h6):(1'h1)]) : $unsigned(reg365[(5'h13):(4'ha)])) : (!reg340[(2'h2):(1'h0)]));
          for (forvar370 = (1'h0); (forvar370 < (1'h0)); forvar370 = (forvar370 + (1'h1)))
            begin
              reg371 <= ((($unsigned($signed(reg367)) <<< reg332[(3'h5):(1'h0)]) > {$signed((reg341 ?
                          (8'ha7) : reg337))}) ?
                  reg303 : reg305[(4'h9):(3'h5)]);
              reg372 <= {reg336,
                  (^~$unsigned(({(8'ha0)} > reg369[(2'h3):(1'h0)])))};
            end
        end
      reg373 <= ((($unsigned(reg321[(4'hf):(3'h4)]) + (reg304[(4'hf):(4'h9)] ?
          $unsigned(reg315) : wire277[(1'h1):(1'h0)])) >> $signed((reg334 > reg305))) - $unsigned((!$signed(wire279[(4'he):(3'h4)]))));
      reg374 <= (reg369[(1'h0):(1'h0)] ?
          ((~|$unsigned($signed(forvar370))) ~^ {({reg357,
                  reg368} <= $unsigned(reg373))}) : reg351[(5'h11):(2'h2)]);
      reg375 <= (^~($unsigned((8'hac)) ?
          $unsigned($signed((reg358 ?
              reg284 : reg345))) : ($unsigned((~|reg367)) | (reg331[(3'h4):(2'h3)] - ((8'h9e) != reg295)))));
    end
  always
    @(posedge clk) begin
      if ($signed((reg303 ?
          $signed({(&reg320), wire279}) : (~(reg358[(1'h1):(1'h0)] ?
              {reg284} : (~reg330))))))
        begin
          reg376 <= reg306;
          for (forvar377 = (1'h0); (forvar377 < (3'h4)); forvar377 = (forvar377 + (1'h1)))
            begin
              reg378 <= $signed(reg295[(1'h1):(1'h0)]);
              reg379 <= (($signed((reg304 ?
                      {(8'h9e)} : $unsigned(reg357))) ^~ wire319) ?
                  reg287[(3'h6):(3'h4)] : $unsigned((((wire280 ?
                          reg337 : (8'hae)) + $unsigned((8'h9f))) ?
                      {(reg305 ? reg304 : reg378)} : reg327)));
            end
          reg380 = (^(reg308 ?
              reg321[(2'h3):(2'h3)] : (($signed(reg374) || reg289[(3'h5):(1'h0)]) >> $unsigned(reg341))));
          reg381 <= $signed((reg375[(1'h1):(1'h1)] | ($unsigned($signed(reg330)) ?
              (8'hb6) : $unsigned((reg378 | wire279)))));
        end
      else
        begin
          reg376 <= ($signed($unsigned((&((8'hbc) ? (8'hb1) : (8'ha3))))) ?
              $signed(reg320[(3'h5):(2'h2)]) : $unsigned($unsigned({{wire279,
                      reg358},
                  {reg371, wire319}})));
          for (forvar377 = (1'h0); (forvar377 < (2'h3)); forvar377 = (forvar377 + (1'h1)))
            begin
              reg380 = {($signed(reg345) ? reg306 : $signed(reg330)),
                  (^~{$signed((reg296 * wire278))})};
              reg381 <= reg305;
            end
        end
      for (forvar382 = (1'h0); (forvar382 < (2'h2)); forvar382 = (forvar382 + (1'h1)))
        begin
          for (forvar383 = (1'h0); (forvar383 < (2'h3)); forvar383 = (forvar383 + (1'h1)))
            begin
              reg384 = (($unsigned($signed(reg285[(2'h2):(1'h1)])) & (^forvar383[(4'h8):(3'h5)])) ?
                  {{$signed((reg379 ? (7'h43) : wire280)), reg345},
                      (~reg340[(2'h2):(1'h1)])} : (reg285 ?
                      $signed(((+reg295) << (reg372 ~^ reg381))) : $unsigned((^{reg369,
                          wire280}))));
            end
          reg385 <= {{{reg306[(3'h5):(2'h2)], $signed((reg297 * reg376))}},
              {(~^$unsigned((8'ha4))), {reg342, {$unsigned(reg341)}}}};
          reg386 = $unsigned((((|(&reg306)) ?
                  reg337[(2'h3):(2'h2)] : ({reg342, wire278} ?
                      (reg351 & reg299) : reg309[(3'h7):(3'h5)])) ?
              reg379 : (&(|(reg354 ? reg305 : reg327)))));
          if (($signed({(reg342 != (8'hb9)), wire280}) ?
              (~|reg284[(4'h8):(2'h3)]) : (reg340[(1'h0):(1'h0)] ?
                  {((reg337 ? reg301 : reg348) ~^ (reg289 ? (7'h42) : reg369)),
                      (+(reg340 >> wire280))} : (((~&reg340) ?
                          (!reg332) : reg378[(4'h8):(3'h7)]) ?
                      ({reg336} ?
                          $signed(reg285) : reg374[(4'hc):(1'h0)]) : {{reg385,
                              wire281},
                          $signed((8'ha2))}))))
            begin
              reg387 <= reg289[(3'h7):(2'h2)];
              reg388 <= $signed((forvar382 << ((!((8'h9d) ?
                  (8'hb9) : reg342)) >> ((reg384 ?
                  reg332 : reg341) >= $unsigned((8'hb4))))));
              reg389 <= reg345;
              reg390 = $signed($unsigned(({((7'h42) <= reg295),
                  reg371} ^ (!((8'hba) ? reg331 : reg330)))));
            end
          else
            begin
              reg387 <= (($unsigned((~&(reg376 << wire281))) ?
                  (reg327 ?
                      ($unsigned(reg296) - (reg336 * reg330)) : (8'hb3)) : (~reg357[(3'h4):(1'h0)])) << reg339[(4'h9):(3'h4)]);
              reg390 = $signed((|(-reg327[(1'h1):(1'h1)])));
            end
        end
    end
  always
    @(posedge clk) begin
      reg391 = $signed($signed({reg330,
          (((8'had) ? reg331 : (8'ha1)) ?
              (reg376 ? reg331 : (7'h44)) : $signed(reg330))}));
      reg392 <= ($signed(reg359) > reg379[(3'h5):(3'h5)]);
      reg393 <= ($unsigned((~|{reg336,
          reg341})) + $unsigned($signed((~&(-(8'haf))))));
    end
  always
    @(posedge clk) begin
      reg394 <= ($signed((8'hb6)) ?
          (8'h9d) : ((+(((8'hbf) ^~ reg314) > {(8'h9f),
              wire278})) ^~ (((^~reg369) ?
                  (reg308 ? (8'ha4) : reg378) : (reg372 + reg379)) ?
              {reg342[(4'hf):(4'ha)], $signed(reg378)} : reg385)));
      for (forvar395 = (1'h0); (forvar395 < (2'h3)); forvar395 = (forvar395 + (1'h1)))
        begin
          reg396 <= (reg295 | (~&$signed(reg358[(2'h3):(1'h0)])));
          reg397 = $signed($signed(reg301[(2'h2):(1'h1)]));
          reg398 <= reg345;
          reg399 = (^~reg358);
        end
      for (forvar400 = (1'h0); (forvar400 < (3'h4)); forvar400 = (forvar400 + (1'h1)))
        begin
          reg401 <= {(~(reg317 ?
                  reg308[(3'h4):(1'h0)] : ((~reg314) ?
                      (^(8'ha2)) : $signed(wire319))))};
          reg402 <= (&(^~reg394));
          reg403 = (8'hbe);
        end
      reg404 = $unsigned(reg342[(4'hb):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg405 <= $unsigned((((|reg358) | ((reg314 << wire279) ^ {reg351})) ?
          {(reg305[(3'h4):(3'h4)] ?
                  $signed(reg285) : ((8'ha0) ?
                      reg345 : reg285))} : reg354[(4'hf):(4'h9)]));
      reg406 <= reg385[(3'h6):(2'h2)];
      reg407 <= (~^(^reg378));
      for (forvar408 = (1'h0); (forvar408 < (3'h4)); forvar408 = (forvar408 + (1'h1)))
        begin
          reg409 <= ((({{reg321, reg355}} ?
                  $signed(reg374[(4'h8):(4'h8)]) : reg369) ^~ ($unsigned(reg367) ?
                  reg372 : $unsigned(reg357))) ?
              {(reg330[(1'h0):(1'h0)] ?
                      ((reg339 + reg372) == wire281[(4'he):(3'h4)]) : (-((8'hb3) ?
                          reg348 : reg324)))} : ($unsigned(reg299[(3'h7):(1'h1)]) ?
                  ((reg284 >= (8'ha2)) ~^ reg340) : $signed(reg334[(4'h9):(2'h2)])));
        end
    end
  always
    @(posedge clk) begin
      reg410 <= reg396;
    end
  always
    @(posedge clk) begin
      reg411 <= $unsigned(($unsigned({(~&reg401)}) <<< {reg306}));
      reg412 <= $signed({(reg284[(1'h0):(1'h0)] ?
              ((^~reg358) - reg314) : (~^$signed(reg299)))});
    end
  always
    @(posedge clk) begin
      for (forvar413 = (1'h0); (forvar413 < (3'h4)); forvar413 = (forvar413 + (1'h1)))
        begin
          reg414 <= (reg388[(1'h0):(1'h0)] ?
              (reg378 >> ({((7'h41) ? (8'hb3) : reg337)} ?
                  $unsigned($unsigned(reg375)) : (reg393 >= $signed(reg330)))) : {(+$signed(reg392))});
        end
      for (forvar415 = (1'h0); (forvar415 < (1'h1)); forvar415 = (forvar415 + (1'h1)))
        begin
          reg416 <= (reg396[(1'h1):(1'h1)] ?
              reg299 : ((8'ha1) ? $signed(reg286) : {reg369[(3'h7):(2'h3)]}));
          reg417 = {$signed(reg285)};
        end
      reg418 <= $unsigned({reg321});
      reg419 <= $signed({reg375[(5'h13):(4'hc)]});
    end
  assign wire420 = reg341;
  always
    @(posedge clk) begin
      for (forvar421 = (1'h0); (forvar421 < (2'h3)); forvar421 = (forvar421 + (1'h1)))
        begin
          reg422 <= (~^(((reg286[(1'h0):(1'h0)] & (reg379 == reg289)) >= (reg367 ?
                  (-reg396) : {(8'ha6)})) ?
              ((wire279 <= (|(8'hbe))) - (8'haa)) : (|reg309)));
          for (forvar423 = (1'h0); (forvar423 < (2'h2)); forvar423 = (forvar423 + (1'h1)))
            begin
              reg424 = $unsigned((8'hae));
            end
          reg425 <= (|((&{{reg357, reg424}, reg365}) > (($unsigned(reg309) ?
              reg292[(4'hf):(2'h3)] : $unsigned(reg372)) << $signed($signed(reg339)))));
          reg426 = $unsigned((reg292[(2'h3):(1'h0)] + $unsigned(reg398)));
          reg427 <= (($unsigned(reg348) ?
              (((reg405 ? reg374 : (8'ha7)) ?
                  {reg287,
                      (8'ha0)} : reg327) < (reg296[(3'h5):(2'h2)] > wire277[(4'ha):(4'ha)])) : ((-(8'ha1)) >= $signed(reg308[(1'h0):(1'h0)]))) ^ ((($signed(reg373) ?
              reg407 : $unsigned(reg378)) > (reg359[(4'ha):(3'h7)] ?
              $signed(forvar421) : $unsigned(wire420))) >>> wire281));
        end
    end
  always
    @(posedge clk) begin
      reg428 <= $unsigned(reg289[(3'h4):(1'h1)]);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module96
#(parameter param272 = (|((((|(8'ha5)) <= {(8'had), (8'hbb)}) ? (^~(!(8'hb6))) : (((7'h41) ~^ (8'hb6)) ? (&(8'hb0)) : ((8'haf) ~^ (7'h40)))) ? (-(((8'ha7) & (8'hb0)) ? ((8'hbe) << (8'h9f)) : (7'h41))) : {(8'ha4)})))
(y, clk, wire101, wire100, wire99, wire98, wire97);
  output wire [(32'h8ce):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hb):(1'h0)] wire101;
  input wire [(4'he):(1'h0)] wire100;
  input wire signed [(5'h12):(1'h0)] wire99;
  input wire signed [(4'hc):(1'h0)] wire98;
  input wire signed [(4'hc):(1'h0)] wire97;
  wire signed [(4'hc):(1'h0)] wire271;
  wire [(3'h7):(1'h0)] wire143;
  reg signed [(3'h5):(1'h0)] reg269 = (1'h0);
  reg [(2'h2):(1'h0)] reg267 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg266 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg263 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg259 = (1'h0);
  reg [(4'hf):(1'h0)] reg258 = (1'h0);
  reg [(4'hf):(1'h0)] reg257 = (1'h0);
  reg [(5'h11):(1'h0)] reg255 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg253 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg251 = (1'h0);
  reg [(5'h15):(1'h0)] reg250 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg247 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg246 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg241 = (1'h0);
  reg [(4'hd):(1'h0)] reg239 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg238 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg235 = (1'h0);
  reg [(5'h15):(1'h0)] reg234 = (1'h0);
  reg [(4'hd):(1'h0)] reg231 = (1'h0);
  reg [(4'hb):(1'h0)] reg227 = (1'h0);
  reg [(5'h12):(1'h0)] reg226 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg224 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg222 = (1'h0);
  reg [(5'h10):(1'h0)] reg219 = (1'h0);
  reg [(2'h2):(1'h0)] reg218 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg215 = (1'h0);
  reg [(3'h7):(1'h0)] reg212 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg210 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg209 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg205 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg198 = (1'h0);
  reg [(5'h15):(1'h0)] reg202 = (1'h0);
  reg [(5'h11):(1'h0)] reg199 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg197 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg193 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg192 = (1'h0);
  reg [(4'ha):(1'h0)] reg191 = (1'h0);
  reg [(3'h5):(1'h0)] reg189 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg185 = (1'h0);
  reg [(5'h13):(1'h0)] reg184 = (1'h0);
  reg [(5'h12):(1'h0)] reg183 = (1'h0);
  reg [(3'h4):(1'h0)] reg182 = (1'h0);
  reg [(5'h13):(1'h0)] reg181 = (1'h0);
  reg [(5'h12):(1'h0)] reg178 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg177 = (1'h0);
  reg [(4'h8):(1'h0)] reg176 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg174 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg173 = (1'h0);
  reg [(5'h14):(1'h0)] reg172 = (1'h0);
  reg [(5'h15):(1'h0)] reg168 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg167 = (1'h0);
  reg [(4'he):(1'h0)] reg166 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg165 = (1'h0);
  reg signed [(4'he):(1'h0)] reg164 = (1'h0);
  reg [(4'h8):(1'h0)] reg162 = (1'h0);
  reg [(3'h6):(1'h0)] reg160 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg159 = (1'h0);
  reg [(4'he):(1'h0)] reg152 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg151 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg150 = (1'h0);
  reg [(3'h6):(1'h0)] reg147 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg146 = (1'h0);
  reg [(4'hd):(1'h0)] reg145 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg144 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg142 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg141 = (1'h0);
  reg [(4'hf):(1'h0)] reg138 = (1'h0);
  reg [(4'h8):(1'h0)] reg136 = (1'h0);
  reg [(4'hc):(1'h0)] reg129 = (1'h0);
  reg [(4'hc):(1'h0)] reg127 = (1'h0);
  reg [(5'h14):(1'h0)] reg126 = (1'h0);
  reg [(3'h5):(1'h0)] reg121 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg125 = (1'h0);
  reg [(5'h15):(1'h0)] reg123 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg120 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg118 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg117 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg116 = (1'h0);
  reg signed [(4'he):(1'h0)] reg115 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg114 = (1'h0);
  reg signed [(4'he):(1'h0)] reg113 = (1'h0);
  reg [(5'h10):(1'h0)] reg111 = (1'h0);
  reg [(5'h12):(1'h0)] reg109 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg108 = (1'h0);
  reg [(3'h6):(1'h0)] reg107 = (1'h0);
  reg [(5'h14):(1'h0)] reg106 = (1'h0);
  reg [(5'h15):(1'h0)] reg102 = (1'h0);
  reg [(5'h12):(1'h0)] reg270 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg268 = (1'h0);
  reg [(4'hb):(1'h0)] reg265 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar264 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar262 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar261 = (1'h0);
  reg [(4'hb):(1'h0)] reg260 = (1'h0);
  reg [(3'h4):(1'h0)] forvar256 = (1'h0);
  reg [(3'h6):(1'h0)] reg254 = (1'h0);
  reg [(4'hd):(1'h0)] forvar252 = (1'h0);
  reg [(4'hb):(1'h0)] reg249 = (1'h0);
  reg [(2'h2):(1'h0)] reg248 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg245 = (1'h0);
  reg [(4'hd):(1'h0)] forvar244 = (1'h0);
  reg [(4'ha):(1'h0)] reg243 = (1'h0);
  reg [(3'h6):(1'h0)] reg242 = (1'h0);
  reg [(4'he):(1'h0)] forvar237 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg237 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg236 = (1'h0);
  reg [(4'ha):(1'h0)] reg233 = (1'h0);
  reg [(4'h9):(1'h0)] reg232 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar230 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg229 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg228 = (1'h0);
  reg [(3'h6):(1'h0)] forvar225 = (1'h0);
  reg [(5'h11):(1'h0)] reg223 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar221 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar220 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar217 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg216 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg214 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg213 = (1'h0);
  reg [(4'hd):(1'h0)] reg211 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg208 = (1'h0);
  reg [(5'h13):(1'h0)] reg207 = (1'h0);
  reg [(5'h11):(1'h0)] reg206 = (1'h0);
  reg signed [(4'he):(1'h0)] reg204 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg203 = (1'h0);
  reg [(4'hd):(1'h0)] forvar201 = (1'h0);
  reg [(2'h2):(1'h0)] reg200 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar198 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg196 = (1'h0);
  reg [(4'ha):(1'h0)] reg195 = (1'h0);
  reg [(5'h12):(1'h0)] reg194 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg190 = (1'h0);
  reg [(2'h3):(1'h0)] forvar188 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar187 = (1'h0);
  reg [(4'hb):(1'h0)] forvar181 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg180 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg175 = (1'h0);
  reg [(4'hb):(1'h0)] reg186 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar180 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg179 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar175 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg171 = (1'h0);
  reg [(4'h8):(1'h0)] reg170 = (1'h0);
  reg [(4'hb):(1'h0)] forvar169 = (1'h0);
  reg [(5'h14):(1'h0)] reg163 = (1'h0);
  reg [(4'he):(1'h0)] reg161 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar158 = (1'h0);
  reg [(3'h5):(1'h0)] forvar157 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg156 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg155 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg154 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg153 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg149 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg148 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar140 = (1'h0);
  reg [(4'ha):(1'h0)] reg139 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg137 = (1'h0);
  reg [(3'h7):(1'h0)] reg135 = (1'h0);
  reg [(5'h12):(1'h0)] reg134 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg133 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg132 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg131 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg130 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar128 = (1'h0);
  reg [(5'h12):(1'h0)] forvar120 = (1'h0);
  reg [(5'h14):(1'h0)] reg124 = (1'h0);
  reg [(5'h10):(1'h0)] reg122 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar121 = (1'h0);
  reg [(4'h9):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar112 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar105 = (1'h0);
  reg [(4'h9):(1'h0)] forvar104 = (1'h0);
  reg [(5'h10):(1'h0)] reg103 = (1'h0);
  assign y = {wire271,
                 wire143,
                 reg269,
                 reg267,
                 reg266,
                 reg263,
                 reg259,
                 reg258,
                 reg257,
                 reg255,
                 reg253,
                 reg251,
                 reg250,
                 reg247,
                 reg246,
                 reg241,
                 reg239,
                 reg238,
                 reg235,
                 reg234,
                 reg231,
                 reg227,
                 reg226,
                 reg224,
                 reg222,
                 reg219,
                 reg218,
                 reg215,
                 reg212,
                 reg210,
                 reg209,
                 reg205,
                 reg198,
                 reg202,
                 reg199,
                 reg197,
                 reg193,
                 reg192,
                 reg191,
                 reg189,
                 reg185,
                 reg184,
                 reg183,
                 reg182,
                 reg181,
                 reg178,
                 reg177,
                 reg176,
                 reg174,
                 reg173,
                 reg172,
                 reg168,
                 reg167,
                 reg166,
                 reg165,
                 reg164,
                 reg162,
                 reg160,
                 reg159,
                 reg152,
                 reg151,
                 reg150,
                 reg147,
                 reg146,
                 reg145,
                 reg144,
                 reg142,
                 reg141,
                 reg138,
                 reg136,
                 reg129,
                 reg127,
                 reg126,
                 reg121,
                 reg125,
                 reg123,
                 reg120,
                 reg118,
                 reg117,
                 reg116,
                 reg115,
                 reg114,
                 reg113,
                 reg111,
                 reg109,
                 reg108,
                 reg107,
                 reg106,
                 reg102,
                 reg270,
                 reg268,
                 reg265,
                 forvar264,
                 forvar262,
                 forvar261,
                 reg260,
                 forvar256,
                 reg254,
                 forvar252,
                 reg249,
                 reg248,
                 reg245,
                 forvar244,
                 reg243,
                 reg242,
                 forvar237,
                 reg240,
                 reg237,
                 reg236,
                 reg233,
                 reg232,
                 forvar230,
                 reg229,
                 reg228,
                 forvar225,
                 reg223,
                 forvar221,
                 forvar220,
                 forvar217,
                 reg216,
                 reg214,
                 reg213,
                 reg211,
                 reg208,
                 reg207,
                 reg206,
                 reg204,
                 reg203,
                 forvar201,
                 reg200,
                 forvar198,
                 reg196,
                 reg195,
                 reg194,
                 reg190,
                 forvar188,
                 forvar187,
                 forvar181,
                 reg180,
                 reg175,
                 reg186,
                 forvar180,
                 reg179,
                 forvar175,
                 reg171,
                 reg170,
                 forvar169,
                 reg163,
                 reg161,
                 forvar158,
                 forvar157,
                 reg156,
                 reg155,
                 reg154,
                 reg153,
                 reg149,
                 reg148,
                 forvar140,
                 reg139,
                 reg137,
                 reg135,
                 reg134,
                 reg133,
                 reg132,
                 reg131,
                 reg130,
                 forvar128,
                 forvar120,
                 reg124,
                 reg122,
                 forvar121,
                 reg119,
                 forvar112,
                 reg110,
                 forvar105,
                 forvar104,
                 reg103,
                 (1'h0)};
  always
    @(posedge clk) begin
      if ($unsigned((8'ha2)))
        begin
          reg102 <= (($unsigned(wire99) ?
                  (~(wire100 >= $unsigned(wire97))) : $signed(((wire99 ?
                      (8'hb1) : wire97) != (!wire97)))) ?
              $signed($unsigned(({(8'hbf),
                  wire98} - (-wire97)))) : $unsigned($signed($signed((wire100 ?
                  wire101 : wire97)))));
        end
      else
        begin
          reg103 = (&(7'h41));
        end
      for (forvar104 = (1'h0); (forvar104 < (2'h2)); forvar104 = (forvar104 + (1'h1)))
        begin
          for (forvar105 = (1'h0); (forvar105 < (3'h4)); forvar105 = (forvar105 + (1'h1)))
            begin
              reg106 <= ((wire98[(4'hb):(4'ha)] ?
                      reg103 : $signed((wire98[(2'h2):(1'h1)] ?
                          (forvar105 & (8'ha4)) : $unsigned(forvar104)))) ?
                  {$signed((-$unsigned(forvar105)))} : wire98);
              reg107 <= (+$unsigned(wire97[(4'hb):(3'h6)]));
              reg108 <= ($unsigned($unsigned((|$unsigned(wire98)))) ?
                  (!$unsigned(reg106)) : $unsigned($unsigned((~&reg107))));
              reg109 <= $signed((+wire99));
              reg110 = $unsigned({wire97});
            end
          reg111 <= $unsigned(((reg108 + forvar104[(3'h6):(3'h4)]) != $unsigned($signed((~^wire98)))));
          for (forvar112 = (1'h0); (forvar112 < (2'h2)); forvar112 = (forvar112 + (1'h1)))
            begin
              reg113 <= ($unsigned({$signed((wire101 ~^ (8'ha4)))}) ?
                  (~&reg103) : ((reg109[(1'h0):(1'h0)] << {reg106[(4'hb):(4'h9)]}) ?
                      (((&reg110) >>> reg109) >> reg111[(4'hd):(3'h6)]) : wire98));
              reg114 <= (8'hb2);
              reg115 <= (8'hb8);
            end
          reg116 <= reg113;
        end
      reg117 <= ((forvar104[(1'h1):(1'h0)] ?
          {({(8'hbe), reg103} ? (wire100 ? reg110 : reg115) : (8'ha5)),
              $unsigned(reg107)} : (~&(~^((8'ha3) == (8'h9d))))) || forvar104[(3'h5):(3'h4)]);
      reg118 <= reg117[(4'hf):(2'h2)];
    end
  always
    @(posedge clk) begin
      reg119 = (reg109 ?
          $unsigned(reg106[(5'h11):(2'h3)]) : wire97[(3'h5):(2'h2)]);
      if (reg113[(3'h7):(2'h2)])
        begin
          reg120 <= $signed(({($signed(reg107) ? wire97 : $unsigned(wire98)),
              $unsigned(reg108)} < $unsigned((reg119 ?
              (reg116 ^ reg115) : (8'ha3)))));
          for (forvar121 = (1'h0); (forvar121 < (2'h2)); forvar121 = (forvar121 + (1'h1)))
            begin
              reg122 = (~(&(^($unsigned(reg117) ?
                  $unsigned((8'hbc)) : reg107))));
              reg123 <= $signed(forvar121[(1'h1):(1'h0)]);
              reg124 = reg106[(1'h0):(1'h0)];
              reg125 <= ((&($unsigned($signed(wire98)) ?
                      {$unsigned(reg122)} : ((reg102 | (7'h43)) ?
                          (7'h43) : reg117))) ?
                  $unsigned((^~(reg124[(4'h8):(1'h1)] << $unsigned(reg114)))) : $unsigned($signed((reg106 - (~reg106)))));
            end
        end
      else
        begin
          for (forvar120 = (1'h0); (forvar120 < (3'h4)); forvar120 = (forvar120 + (1'h1)))
            begin
              reg121 <= $signed($unsigned($unsigned({(8'h9c)})));
              reg123 <= (|$unsigned($signed(reg107)));
              reg125 <= (+($unsigned(($unsigned(reg119) & reg114[(1'h0):(1'h0)])) ?
                  ($unsigned((~&reg113)) ?
                      reg118[(1'h0):(1'h0)] : reg123) : ((~(reg125 ?
                      reg115 : wire98)) | reg114[(2'h3):(2'h2)])));
              reg126 <= (^(7'h44));
              reg127 <= reg118;
            end
          for (forvar128 = (1'h0); (forvar128 < (3'h4)); forvar128 = (forvar128 + (1'h1)))
            begin
              reg129 <= (^~reg123);
              reg130 = ($unsigned($unsigned(((reg124 - reg120) ?
                      $signed(reg111) : (!reg122)))) ?
                  reg116 : {(~&reg102[(4'hc):(1'h0)]), reg121});
              reg131 = $signed($unsigned(($unsigned((reg107 <<< (7'h41))) ?
                  ((reg121 ?
                      reg115 : reg124) ^ forvar128[(4'hc):(1'h0)]) : forvar120[(1'h1):(1'h1)])));
              reg132 = (($unsigned(((reg115 <= forvar121) ?
                          reg125[(4'h8):(3'h7)] : reg126)) ?
                      (reg125[(1'h1):(1'h1)] - reg113[(3'h6):(3'h4)]) : reg125) ?
                  {(|(((8'hbf) ?
                          wire100 : forvar128) != (wire99 + reg102)))} : $unsigned((($signed(reg116) ?
                          (~^reg131) : (8'hb0)) ?
                      $signed((reg124 ?
                          reg114 : reg111)) : $signed(reg126[(3'h6):(3'h6)]))));
              reg133 = reg102[(4'hf):(4'hd)];
            end
          reg134 = $unsigned($signed(reg109[(4'h9):(4'h8)]));
          reg135 = $unsigned($signed((reg107[(2'h2):(1'h1)] ?
              (~|$signed(reg115)) : reg115)));
        end
      if ((reg120 ?
          $unsigned(((~^(~reg132)) << {reg133[(1'h1):(1'h0)],
              ((8'hb2) ?
                  reg125 : wire100)})) : ({reg123} <= reg111[(2'h3):(1'h0)])))
        begin
          reg136 <= $signed((!$signed((~^(~|(8'haf))))));
          reg137 = (reg102[(3'h6):(3'h6)] ?
              reg125 : (+{($signed(wire99) > (reg106 ? (8'hb1) : reg106))}));
        end
      else
        begin
          reg136 <= (-(reg111[(4'hd):(4'ha)] ?
              ($unsigned((reg102 ?
                  reg117 : reg106)) >= {reg126}) : $signed(reg116)));
          reg137 = (reg106[(4'hc):(4'h8)] ?
              {$signed((^~(reg118 & reg111))),
                  (+(reg109 ?
                      (wire99 > reg135) : $unsigned(reg130)))} : ({reg113} != reg108));
          reg138 <= (+reg126[(4'ha):(3'h5)]);
        end
      reg139 = reg109;
    end
  always
    @(posedge clk) begin
      for (forvar140 = (1'h0); (forvar140 < (2'h2)); forvar140 = (forvar140 + (1'h1)))
        begin
          reg141 <= (((!($signed(reg136) ?
                  $unsigned(reg138) : reg118[(1'h1):(1'h0)])) + $unsigned((reg106[(5'h13):(4'ha)] != (reg120 >> reg138)))) ?
              $unsigned({((-reg120) ? wire97 : (&(8'hbc))),
                  (-$signed(reg123))}) : ((reg116[(3'h7):(1'h0)] ?
                      {$signed(reg121)} : {{reg121, reg107}}) ?
                  $unsigned(reg114[(1'h0):(1'h0)]) : ({$signed((8'hb6))} * ($unsigned(reg117) ?
                      (reg120 - reg127) : $unsigned((8'hb5))))));
        end
      reg142 <= $signed((reg111[(4'ha):(2'h2)] << (reg109 ?
          ($unsigned(reg116) ?
              reg118[(2'h3):(1'h0)] : reg123[(5'h14):(5'h13)]) : (-(reg107 & reg121)))));
    end
  assign wire143 = $unsigned(reg116[(3'h5):(2'h2)]);
  always
    @(posedge clk) begin
      reg144 <= ($signed(reg125[(2'h2):(2'h2)]) ?
          reg138[(2'h3):(1'h0)] : reg114[(1'h1):(1'h1)]);
      if (((~&$signed((|reg102[(5'h11):(4'he)]))) && (({(reg108 ^ (8'ha6)),
              (+reg116)} != (reg129 ?
              reg108[(4'ha):(3'h4)] : (wire97 & reg127))) ?
          (~&reg109) : $unsigned((reg116 ? (&reg121) : (^wire101))))))
        begin
          reg145 <= ((reg111[(5'h10):(3'h7)] | ($signed({reg109}) ?
              $unsigned(wire100[(3'h6):(1'h0)]) : $unsigned(reg114))) + (reg115 ?
              ($signed($signed(reg129)) > $signed($signed(reg116))) : (~&reg118)));
        end
      else
        begin
          reg145 <= (!(&reg111[(4'hf):(3'h6)]));
          if (reg107)
            begin
              reg146 <= ((-reg109) + $unsigned(reg113[(1'h0):(1'h0)]));
            end
          else
            begin
              reg146 <= reg145;
              reg147 <= $signed($unsigned($unsigned(reg126[(3'h4):(2'h2)])));
            end
        end
      if ((!((reg113 + $signed((reg116 ?
          reg107 : reg113))) ~^ ($signed(wire97[(4'h9):(2'h2)]) ?
          ((~|reg109) ?
              $unsigned(reg111) : $unsigned(reg106)) : (^~$unsigned(reg113))))))
        begin
          reg148 = ($signed({(~&reg113[(2'h2):(2'h2)]),
              reg106[(4'hb):(3'h5)]}) | (+(!($signed(reg117) ?
              (reg141 ^~ reg121) : (wire143 != (8'ha6))))));
          if ($signed({(+((~|reg145) >= reg121[(1'h0):(1'h0)]))}))
            begin
              reg149 = (($unsigned(wire99) >= (~|(~^$signed(wire143)))) && (~|wire100[(4'h9):(3'h4)]));
              reg150 <= (~{((8'hb6) || reg146[(3'h7):(3'h5)]), reg109});
              reg151 <= $signed($signed(reg114[(1'h0):(1'h0)]));
              reg152 <= wire143[(2'h3):(2'h3)];
            end
          else
            begin
              reg150 <= (($signed(reg136[(3'h5):(1'h1)]) + ($signed($unsigned(reg144)) ?
                  $unsigned({reg118}) : reg123[(3'h7):(3'h5)])) >= (~|$unsigned((((7'h44) >>> wire101) ?
                  reg107 : $signed(wire100)))));
              reg153 = $signed(($signed(reg144) != reg129));
              reg154 = (-reg127[(2'h2):(1'h0)]);
              reg155 = reg147;
              reg156 = (^~wire97);
            end
        end
      else
        begin
          reg148 = ($unsigned($signed(wire98)) ?
              ((reg146 != (^~reg106[(3'h6):(1'h0)])) >> reg146) : (|(|$signed(reg152))));
        end
      for (forvar157 = (1'h0); (forvar157 < (1'h0)); forvar157 = (forvar157 + (1'h1)))
        begin
          for (forvar158 = (1'h0); (forvar158 < (2'h3)); forvar158 = (forvar158 + (1'h1)))
            begin
              reg159 <= reg108[(4'hc):(3'h4)];
              reg160 <= $signed((|reg136[(3'h5):(3'h5)]));
            end
          reg161 = (~^$unsigned(($unsigned((wire97 > reg153)) ?
              (8'ha6) : ($unsigned(reg118) ?
                  (^(8'hbd)) : (reg154 ? reg109 : (8'ha5))))));
          if (($unsigned((-reg129)) <<< reg151[(4'h8):(3'h6)]))
            begin
              reg162 <= $signed($signed($signed(reg149[(1'h1):(1'h1)])));
            end
          else
            begin
              reg162 <= (&({((wire101 ? reg146 : reg109) ?
                          $unsigned((8'hb4)) : $signed(wire101)),
                      wire98} ?
                  (|(~|$signed((8'h9e)))) : $unsigned(({reg161, reg145} ?
                      (^~reg155) : (wire100 * reg154)))));
              reg163 = reg120;
              reg164 <= $signed(((reg111 ^ $signed((reg102 ?
                      (8'h9d) : reg138))) ?
                  $signed(reg149[(1'h0):(1'h0)]) : (-reg152[(1'h1):(1'h0)])));
              reg165 <= $unsigned($signed({(^~(wire101 & reg155))}));
              reg166 <= (|$signed(reg138[(4'hc):(1'h0)]));
            end
          reg167 <= ($unsigned((reg149[(2'h3):(1'h1)] << $unsigned(reg141))) ?
              $unsigned((((~^reg156) | (reg152 ? reg156 : reg109)) ?
                  ((reg144 ? reg129 : reg164) ?
                      reg160[(2'h3):(1'h0)] : $unsigned(reg113)) : reg109[(5'h12):(5'h10)])) : reg129);
          reg168 <= (reg121[(3'h5):(2'h3)] + $signed(forvar157));
        end
    end
  always
    @(posedge clk) begin
      if (reg120)
        begin
          for (forvar169 = (1'h0); (forvar169 < (2'h2)); forvar169 = (forvar169 + (1'h1)))
            begin
              reg170 = (reg142 ? reg142[(4'hb):(2'h3)] : reg106[(4'hc):(2'h3)]);
              reg171 = $signed(reg166);
              reg172 <= reg123[(1'h1):(1'h0)];
              reg173 <= $unsigned(reg120);
              reg174 <= $signed((+reg165[(2'h3):(2'h3)]));
            end
          for (forvar175 = (1'h0); (forvar175 < (1'h0)); forvar175 = (forvar175 + (1'h1)))
            begin
              reg176 <= (^~$unsigned(reg167));
              reg177 <= reg168[(2'h2):(2'h2)];
              reg178 <= reg168;
              reg179 = reg170[(3'h6):(3'h4)];
            end
          for (forvar180 = (1'h0); (forvar180 < (2'h2)); forvar180 = (forvar180 + (1'h1)))
            begin
              reg181 <= (8'ha1);
              reg182 <= ((~^$signed(reg146[(4'hb):(2'h3)])) ?
                  (-(|($unsigned(forvar180) ?
                      reg167[(3'h5):(2'h2)] : reg167))) : reg166[(1'h1):(1'h1)]);
              reg183 <= wire99;
              reg184 <= (wire100[(2'h3):(2'h2)] <= ((-$signed($signed(reg171))) ?
                  ($signed(forvar175[(3'h6):(2'h2)]) >= forvar180[(2'h3):(2'h3)]) : (-reg182)));
            end
          reg185 <= ($signed(reg159) ? (^reg116) : $unsigned((^~(~|{reg142}))));
          reg186 = reg142[(4'hd):(4'h8)];
        end
      else
        begin
          for (forvar169 = (1'h0); (forvar169 < (2'h3)); forvar169 = (forvar169 + (1'h1)))
            begin
              reg172 <= (~&(wire99 >= (reg111 ? $signed({(8'h9e)}) : reg184)));
              reg173 <= reg159;
              reg175 = ($unsigned({$signed(((8'had) ? reg150 : reg179))}) ?
                  $signed($unsigned((reg173 ^~ (forvar180 > forvar169)))) : $signed(((7'h41) ?
                      reg136[(1'h1):(1'h0)] : $signed($signed(reg146)))));
              reg176 <= (($signed(((|reg173) != $unsigned(reg114))) ?
                  $unsigned(($signed(reg129) < wire97)) : (^$unsigned(reg146[(1'h0):(1'h0)]))) & (reg168[(4'hc):(3'h5)] ?
                  $unsigned((reg160 + (reg127 ? reg123 : wire99))) : (((7'h43) ?
                          (reg166 ? (8'h9e) : reg127) : (reg107 >= (8'hae))) ?
                      $unsigned((forvar175 ?
                          reg164 : reg127)) : (reg109[(5'h12):(4'hd)] ?
                          (^~reg109) : (reg167 ? reg117 : (8'ha1))))));
              reg177 <= reg184[(3'h5):(2'h3)];
            end
          reg179 = $signed(reg129);
          reg180 = reg108[(4'h8):(2'h3)];
          for (forvar181 = (1'h0); (forvar181 < (3'h4)); forvar181 = (forvar181 + (1'h1)))
            begin
              reg182 <= $unsigned($unsigned($unsigned(((~^(7'h44)) <<< {wire98,
                  forvar169}))));
              reg186 = (((~|{$unsigned(reg159)}) ?
                  (~$unsigned(forvar175[(4'h9):(4'h8)])) : reg177[(4'h8):(3'h5)]) ^ $unsigned((reg136 ?
                  reg126 : (wire101[(3'h7):(1'h0)] ^ (reg102 - reg127)))));
            end
        end
      for (forvar187 = (1'h0); (forvar187 < (1'h0)); forvar187 = (forvar187 + (1'h1)))
        begin
          for (forvar188 = (1'h0); (forvar188 < (1'h0)); forvar188 = (forvar188 + (1'h1)))
            begin
              reg189 <= reg175[(2'h3):(2'h3)];
            end
        end
      reg190 = ({reg174} >>> (8'ha2));
      reg191 <= ($unsigned(reg141) >= reg117[(4'hb):(4'h8)]);
    end
  always
    @(posedge clk) begin
      reg192 <= reg117;
      reg193 <= $signed((({reg114} ?
              ((~|reg189) ?
                  (reg127 ~^ reg152) : (|(7'h40))) : $unsigned($signed((8'hb6)))) ?
          $signed(reg183[(3'h4):(1'h0)]) : wire97));
      reg194 = reg106[(1'h0):(1'h0)];
      reg195 = reg106[(2'h2):(1'h0)];
    end
  always
    @(posedge clk) begin
      reg196 = $signed($signed(((reg181 || (|(8'ha2))) ?
          $unsigned(reg184[(4'hc):(4'h9)]) : $unsigned($unsigned(reg117)))));
    end
  always
    @(posedge clk) begin
      if ($unsigned(reg126[(4'hf):(3'h6)]))
        begin
          reg197 <= (~|(reg160 ? reg109 : (|((!reg172) << $signed(reg166)))));
          for (forvar198 = (1'h0); (forvar198 < (1'h0)); forvar198 = (forvar198 + (1'h1)))
            begin
              reg199 <= {(&reg177[(1'h0):(1'h0)]), (8'h9e)};
              reg200 = {{((~&reg181[(4'hd):(1'h0)]) ~^ {$unsigned(reg116),
                          (~^wire100)}),
                      (reg174 ? reg142 : $unsigned({reg127}))},
                  forvar198};
            end
          for (forvar201 = (1'h0); (forvar201 < (1'h0)); forvar201 = (forvar201 + (1'h1)))
            begin
              reg202 <= $signed($unsigned((-((reg108 && reg151) ^ (reg165 ?
                  (8'hb1) : (8'h9d))))));
              reg203 = $unsigned(reg185[(5'h10):(4'h9)]);
              reg204 = reg159[(1'h1):(1'h1)];
            end
        end
      else
        begin
          reg197 <= reg204[(3'h5):(3'h5)];
          reg198 <= wire101;
          reg200 = (reg123[(4'hd):(4'hc)] <<< (((forvar201[(1'h1):(1'h1)] ?
                  reg164 : (reg118 ? reg198 : reg165)) >> $unsigned({reg126,
                  forvar198})) ?
              $unsigned(((^reg164) ^~ $signed(wire100))) : reg183));
          for (forvar201 = (1'h0); (forvar201 < (2'h3)); forvar201 = (forvar201 + (1'h1)))
            begin
              reg203 = reg147;
              reg205 <= $signed((($signed({reg109,
                  reg202}) < $signed((!reg121))) & reg173[(4'h8):(1'h0)]));
              reg206 = reg151[(4'hd):(4'ha)];
              reg207 = ((|{(reg174 >>> $signed(reg109))}) ^ $unsigned((^reg152[(2'h2):(1'h0)])));
              reg208 = reg123;
            end
          reg209 <= ((wire99 ^~ (-(reg203[(1'h1):(1'h0)] ?
                  reg108 : $signed(reg117)))) ?
              $signed($signed(forvar201)) : ($signed(((reg197 < reg108) ?
                      (!reg160) : $unsigned(reg174))) ?
                  reg204[(2'h3):(1'h1)] : reg126[(5'h10):(4'hb)]));
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned((&$unsigned((~reg172[(5'h11):(4'he)])))))
        begin
          if (((8'hb4) ? reg192[(4'hc):(4'ha)] : reg197[(1'h1):(1'h1)]))
            begin
              reg210 <= reg129;
              reg211 = ({{reg182},
                      (reg210[(2'h3):(1'h0)] < $signed(reg117[(4'hc):(2'h2)]))} ?
                  $signed(reg162) : reg109[(2'h2):(1'h0)]);
              reg212 <= (reg129[(4'ha):(3'h5)] - $signed($signed((reg211 ?
                  $unsigned(reg121) : {reg123}))));
              reg213 = reg168;
              reg214 = (reg211[(4'hb):(4'h9)] == {reg145[(2'h2):(2'h2)],
                  $unsigned((+(8'hb1)))});
            end
          else
            begin
              reg211 = reg121[(3'h4):(3'h4)];
              reg213 = reg212[(1'h0):(1'h0)];
            end
          reg215 <= $signed((~^$signed(((reg109 + reg115) * reg106))));
          reg216 = (reg102[(4'hd):(4'ha)] != $signed($signed(((+reg160) >> (reg121 != (8'hb0))))));
        end
      else
        begin
          reg210 <= wire101;
        end
      for (forvar217 = (1'h0); (forvar217 < (2'h3)); forvar217 = (forvar217 + (1'h1)))
        begin
          reg218 <= ({(-reg145)} ^ reg126[(2'h2):(1'h1)]);
        end
      reg219 <= reg182;
      for (forvar220 = (1'h0); (forvar220 < (2'h2)); forvar220 = (forvar220 + (1'h1)))
        begin
          for (forvar221 = (1'h0); (forvar221 < (2'h2)); forvar221 = (forvar221 + (1'h1)))
            begin
              reg222 <= ((8'hbf) * (~wire98));
              reg223 = reg120;
              reg224 <= $signed(((^~$unsigned((reg184 ?
                  (8'h9c) : (8'hbf)))) << reg125));
            end
          for (forvar225 = (1'h0); (forvar225 < (2'h2)); forvar225 = (forvar225 + (1'h1)))
            begin
              reg226 <= $signed(reg118[(1'h1):(1'h1)]);
              reg227 <= ({$signed({$signed(reg116),
                      reg152[(4'ha):(2'h2)]})} + $unsigned((^~reg107)));
              reg228 = $signed((~^(^reg176[(3'h7):(3'h4)])));
              reg229 = ($unsigned($signed(wire100)) && $signed(reg177));
            end
          for (forvar230 = (1'h0); (forvar230 < (1'h0)); forvar230 = (forvar230 + (1'h1)))
            begin
              reg231 <= (^~$unsigned($unsigned(reg167[(1'h1):(1'h0)])));
              reg232 = $unsigned((!$signed(reg181[(4'h9):(2'h3)])));
              reg233 = {$unsigned(reg185[(4'hf):(4'hc)])};
              reg234 <= (reg106[(3'h6):(3'h4)] ?
                  (reg159[(2'h3):(2'h3)] ?
                      (^~$signed($signed(reg147))) : reg107[(2'h2):(1'h0)]) : $unsigned(reg214));
              reg235 <= $unsigned($unsigned($signed($signed($unsigned(reg114)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg236 = ((reg167[(3'h5):(3'h4)] ?
              reg152 : (~&($signed(reg127) == reg199[(1'h0):(1'h0)]))) ?
          reg125[(2'h2):(1'h1)] : {((^~(reg118 ? reg106 : (8'ha6))) ?
                  $signed($signed(reg198)) : (+$unsigned((8'ha0)))),
              $signed($signed(reg174))});
      if (({{reg189[(2'h2):(1'h1)], reg160}} - reg224[(4'hd):(4'ha)]))
        begin
          reg237 = reg236;
          reg238 <= (((~^($unsigned(reg218) ?
                  $signed((8'hac)) : (-reg165))) * (~reg162)) ?
              reg136[(3'h5):(2'h3)] : $unsigned({{(reg174 ? reg176 : reg183),
                      {reg193, reg219}}}));
          if (wire97)
            begin
              reg239 <= {$signed((~^reg142[(4'hd):(4'h9)]))};
            end
          else
            begin
              reg239 <= {reg123};
            end
          reg240 = (($unsigned($signed((^reg191))) ?
              reg167[(3'h4):(2'h3)] : reg102[(4'h8):(3'h6)]) < $signed(($unsigned($unsigned(reg150)) ?
              ({reg136, reg168} ?
                  {reg238, (8'hb1)} : {reg118, reg212}) : ((~(8'ha5)) ?
                  (reg152 >>> reg107) : $signed(wire143)))));
          reg241 <= $signed((~reg165));
        end
      else
        begin
          for (forvar237 = (1'h0); (forvar237 < (3'h4)); forvar237 = (forvar237 + (1'h1)))
            begin
              reg238 <= $signed(((($signed(reg151) || $signed(reg145)) * (8'hb2)) >= reg235[(2'h3):(1'h1)]));
              reg240 = (&$unsigned((reg215 < $signed(reg150[(1'h0):(1'h0)]))));
              reg241 <= $signed($unsigned((~&{$unsigned(reg144)})));
              reg242 = reg152[(4'he):(4'h9)];
              reg243 = reg129[(4'hc):(4'ha)];
            end
          for (forvar244 = (1'h0); (forvar244 < (2'h3)); forvar244 = (forvar244 + (1'h1)))
            begin
              reg245 = $signed(reg120[(4'h9):(2'h3)]);
              reg246 <= $signed(reg106);
              reg247 <= $signed(reg237[(1'h0):(1'h0)]);
              reg248 = reg127[(4'hc):(2'h3)];
              reg249 = (&reg136);
            end
        end
      reg250 <= (~|reg212[(2'h2):(1'h1)]);
    end
  always
    @(posedge clk) begin
      reg251 <= reg106;
      for (forvar252 = (1'h0); (forvar252 < (2'h2)); forvar252 = (forvar252 + (1'h1)))
        begin
          reg253 <= {((((reg162 >= reg151) >= (-(8'hac))) | reg215) ?
                  {reg174,
                      ($unsigned(reg116) ?
                          (reg224 ?
                              reg199 : wire98) : wire97)} : (^{((8'hb9) & reg239)}))};
          reg254 = $unsigned((^~$signed({(reg238 ? wire98 : reg241),
              (reg165 ? reg108 : reg176)})));
          reg255 <= ((reg107 ?
              forvar252[(4'hd):(3'h6)] : (reg210 ?
                  (-$unsigned((8'had))) : reg202)) >> (~&reg168));
        end
      for (forvar256 = (1'h0); (forvar256 < (1'h0)); forvar256 = (forvar256 + (1'h1)))
        begin
          reg257 <= reg106[(3'h5):(2'h2)];
          reg258 <= ((~^$signed(reg239[(4'h8):(4'h8)])) >= ((|(|(&reg123))) ?
              $signed((|(^reg182))) : (reg250 > {$unsigned(reg113),
                  (wire99 ? reg121 : (8'hbc))})));
        end
      reg259 <= {$unsigned(({reg136[(3'h5):(3'h4)],
              (reg254 ? reg126 : (8'hbb))} < $unsigned(reg197[(1'h1):(1'h1)]))),
          (reg113 ? {(~|(&(8'hb8)))} : reg202[(4'hf):(3'h4)])};
    end
  always
    @(posedge clk) begin
      reg260 = reg257;
    end
  always
    @(posedge clk) begin
      for (forvar261 = (1'h0); (forvar261 < (1'h0)); forvar261 = (forvar261 + (1'h1)))
        begin
          for (forvar262 = (1'h0); (forvar262 < (1'h0)); forvar262 = (forvar262 + (1'h1)))
            begin
              reg263 <= (|$signed((8'had)));
            end
          for (forvar264 = (1'h0); (forvar264 < (3'h4)); forvar264 = (forvar264 + (1'h1)))
            begin
              reg265 = ((reg202 ?
                  ((|(~&reg172)) ?
                      $signed((reg108 ? reg108 : reg224)) : {reg165,
                          (reg173 ?
                              reg117 : reg234)}) : ((reg238[(1'h1):(1'h0)] ~^ $signed(forvar262)) ~^ ((reg166 ?
                          reg250 : reg227) ?
                      $unsigned(reg174) : reg246[(2'h3):(1'h1)]))) <<< ($signed(reg197[(1'h1):(1'h1)]) > ((reg235[(3'h7):(2'h2)] >>> $unsigned(reg199)) ?
                  $unsigned($signed(reg146)) : ((reg226 ?
                      reg151 : reg125) > ((8'hbb) ? reg246 : wire100)))));
              reg266 <= reg259[(1'h1):(1'h1)];
            end
          reg267 <= (8'ha6);
          reg268 = (((reg114[(2'h2):(1'h1)] | $unsigned((|reg193))) ^~ ((((8'hbe) < reg257) & reg238) ?
                  $signed((+(8'h9e))) : reg176)) ?
              (8'hb3) : reg159);
        end
      reg269 <= reg162;
      reg270 = $signed({wire100});
    end
  assign wire271 = $signed({(~(reg116 ?
                           reg191[(3'h6):(2'h2)] : $signed(reg267)))});
endmodule