(* use_dsp48="no" *) (* use_dsp="no" *) module top
#(parameter param1393 = (((~|(~(^~(8'had)))) >>> (^~((~(8'hab)) ? (!(8'haa)) : (~(8'ha8))))) < (((((8'ha3) * (8'hbb)) ? (~(8'had)) : (8'hb5)) ? (~&{(8'hac), (8'hb9)}) : (((7'h45) ? (7'h44) : (8'ha3)) ? ((8'ha3) ~^ (8'ha2)) : ((7'h40) >> (7'h46)))) + {{(!(7'h49))}})))
(y, clk, wire3, wire2, wire1, wire0);
  output wire [(32'hf99):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h10):(1'h0)] wire3;
  input wire signed [(5'h18):(1'h0)] wire2;
  input wire [(5'h14):(1'h0)] wire1;
  input wire [(5'h15):(1'h0)] wire0;
  wire signed [(5'h14):(1'h0)] wire1389;
  wire signed [(4'hc):(1'h0)] wire1388;
  wire signed [(3'h5):(1'h0)] wire1342;
  wire [(4'hb):(1'h0)] wire1336;
  wire signed [(4'h8):(1'h0)] wire1335;
  wire signed [(4'hb):(1'h0)] wire1291;
  wire [(3'h6):(1'h0)] wire1290;
  wire [(5'h18):(1'h0)] wire1261;
  wire signed [(5'h12):(1'h0)] wire1260;
  wire [(5'h17):(1'h0)] wire1211;
  wire [(5'h10):(1'h0)] wire120;
  wire [(4'hc):(1'h0)] wire4;
  reg [(2'h3):(1'h0)] reg1392 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1387 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1384 = (1'h0);
  reg [(5'h13):(1'h0)] reg1382 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1379 = (1'h0);
  reg [(5'h17):(1'h0)] reg1378 = (1'h0);
  reg [(4'hb):(1'h0)] reg1376 = (1'h0);
  reg [(5'h18):(1'h0)] reg1375 = (1'h0);
  reg [(4'hc):(1'h0)] reg1374 = (1'h0);
  reg [(5'h11):(1'h0)] reg1372 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1370 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1368 = (1'h0);
  reg [(5'h16):(1'h0)] reg1365 = (1'h0);
  reg [(4'hb):(1'h0)] reg1356 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1355 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1354 = (1'h0);
  reg [(4'he):(1'h0)] reg1351 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1350 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1348 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1347 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1344 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1341 = (1'h0);
  reg [(4'hc):(1'h0)] reg1337 = (1'h0);
  reg [(3'h5):(1'h0)] reg1334 = (1'h0);
  reg [(5'h14):(1'h0)] reg1332 = (1'h0);
  reg [(2'h2):(1'h0)] reg1331 = (1'h0);
  reg [(3'h5):(1'h0)] reg1330 = (1'h0);
  reg [(5'h10):(1'h0)] reg1327 = (1'h0);
  reg [(4'h9):(1'h0)] reg1323 = (1'h0);
  reg [(5'h17):(1'h0)] reg1321 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1320 = (1'h0);
  reg [(3'h4):(1'h0)] reg1314 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1311 = (1'h0);
  reg [(4'hd):(1'h0)] reg1307 = (1'h0);
  reg [(4'he):(1'h0)] reg1306 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1305 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1303 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1300 = (1'h0);
  reg [(5'h17):(1'h0)] reg1296 = (1'h0);
  reg [(4'hc):(1'h0)] reg1295 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1292 = (1'h0);
  reg [(3'h4):(1'h0)] reg1286 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1281 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1278 = (1'h0);
  reg [(5'h10):(1'h0)] reg1277 = (1'h0);
  reg [(4'hd):(1'h0)] reg1276 = (1'h0);
  reg [(5'h16):(1'h0)] reg1274 = (1'h0);
  reg [(4'ha):(1'h0)] reg1271 = (1'h0);
  reg [(4'hc):(1'h0)] reg1269 = (1'h0);
  reg [(3'h6):(1'h0)] reg1267 = (1'h0);
  reg [(4'hc):(1'h0)] reg1266 = (1'h0);
  reg [(3'h4):(1'h0)] reg1263 = (1'h0);
  reg [(3'h6):(1'h0)] reg1259 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1255 = (1'h0);
  reg [(3'h6):(1'h0)] reg1254 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1246 = (1'h0);
  reg [(5'h11):(1'h0)] reg1245 = (1'h0);
  reg [(4'hb):(1'h0)] reg1242 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1240 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1235 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1234 = (1'h0);
  reg [(3'h4):(1'h0)] reg1233 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1229 = (1'h0);
  reg [(3'h5):(1'h0)] reg1228 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1227 = (1'h0);
  reg [(4'h9):(1'h0)] reg1225 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1224 = (1'h0);
  reg [(5'h16):(1'h0)] reg1223 = (1'h0);
  reg [(2'h3):(1'h0)] reg1222 = (1'h0);
  reg [(4'h9):(1'h0)] reg1221 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1216 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1213 = (1'h0);
  reg [(4'h8):(1'h0)] reg116 = (1'h0);
  reg [(2'h3):(1'h0)] reg111 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg110 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg109 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg108 = (1'h0);
  reg [(4'hf):(1'h0)] reg105 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg104 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg101 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg100 = (1'h0);
  reg [(4'h9):(1'h0)] reg99 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg97 = (1'h0);
  reg [(5'h12):(1'h0)] reg95 = (1'h0);
  reg signed [(4'he):(1'h0)] reg93 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg92 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg85 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg91 = (1'h0);
  reg signed [(4'he):(1'h0)] reg89 = (1'h0);
  reg [(5'h10):(1'h0)] reg87 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg83 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg82 = (1'h0);
  reg [(4'h8):(1'h0)] reg81 = (1'h0);
  reg [(4'h9):(1'h0)] reg78 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg75 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg74 = (1'h0);
  reg [(5'h14):(1'h0)] reg72 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg70 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg69 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg67 = (1'h0);
  reg [(4'hd):(1'h0)] reg63 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg57 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg55 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg49 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg45 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg44 = (1'h0);
  reg [(4'hd):(1'h0)] reg43 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg42 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg41 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg40 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg37 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg34 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg31 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg27 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg26 = (1'h0);
  reg [(3'h5):(1'h0)] reg22 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg21 = (1'h0);
  reg [(3'h4):(1'h0)] reg17 = (1'h0);
  reg [(5'h16):(1'h0)] reg16 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg15 = (1'h0);
  reg [(5'h18):(1'h0)] reg14 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg13 = (1'h0);
  reg [(5'h17):(1'h0)] reg11 = (1'h0);
  reg [(4'hb):(1'h0)] reg1391 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1390 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1386 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar1385 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1373 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1368 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1383 = (1'h0);
  reg [(4'he):(1'h0)] reg1381 = (1'h0);
  reg [(4'hd):(1'h0)] reg1380 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1377 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1373 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1371 = (1'h0);
  reg [(5'h16):(1'h0)] reg1369 = (1'h0);
  reg [(4'h9):(1'h0)] reg1367 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1366 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1364 = (1'h0);
  reg [(4'h8):(1'h0)] reg1363 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1362 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1361 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1360 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1359 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1358 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1357 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1354 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1352 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1353 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1352 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1349 = (1'h0);
  reg [(4'hb):(1'h0)] reg1343 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1346 = (1'h0);
  reg [(2'h3):(1'h0)] reg1345 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1343 = (1'h0);
  reg [(2'h3):(1'h0)] reg1340 = (1'h0);
  reg [(3'h4):(1'h0)] reg1339 = (1'h0);
  reg [(4'hd):(1'h0)] reg1338 = (1'h0);
  reg [(4'hd):(1'h0)] reg1333 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1329 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1328 = (1'h0);
  reg [(4'hf):(1'h0)] reg1326 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1325 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1324 = (1'h0);
  reg [(3'h7):(1'h0)] reg1322 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1319 = (1'h0);
  reg [(4'hf):(1'h0)] reg1318 = (1'h0);
  reg [(4'h8):(1'h0)] reg1317 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1316 = (1'h0);
  reg [(4'ha):(1'h0)] reg1315 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1313 = (1'h0);
  reg [(2'h2):(1'h0)] reg1312 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1310 = (1'h0);
  reg [(4'hf):(1'h0)] reg1309 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1308 = (1'h0);
  reg [(5'h16):(1'h0)] reg1304 = (1'h0);
  reg [(5'h13):(1'h0)] reg1302 = (1'h0);
  reg [(5'h18):(1'h0)] reg1301 = (1'h0);
  reg [(3'h6):(1'h0)] reg1299 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1298 = (1'h0);
  reg [(5'h13):(1'h0)] reg1293 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar1292 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1297 = (1'h0);
  reg [(4'h8):(1'h0)] reg1294 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1293 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1289 = (1'h0);
  reg [(3'h7):(1'h0)] reg1288 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1287 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1285 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1284 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1283 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar1282 = (1'h0);
  reg [(4'hc):(1'h0)] reg1280 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1279 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1275 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1273 = (1'h0);
  reg [(3'h7):(1'h0)] reg1272 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1270 = (1'h0);
  reg [(3'h7):(1'h0)] forvar1268 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1265 = (1'h0);
  reg [(5'h15):(1'h0)] reg1264 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1262 = (1'h0);
  reg [(4'hd):(1'h0)] reg1258 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1257 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1256 = (1'h0);
  reg [(5'h12):(1'h0)] forvar1253 = (1'h0);
  reg [(4'hf):(1'h0)] reg1252 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1251 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1250 = (1'h0);
  reg [(4'hb):(1'h0)] forvar1249 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1248 = (1'h0);
  reg [(5'h11):(1'h0)] reg1247 = (1'h0);
  reg [(5'h15):(1'h0)] reg1244 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1243 = (1'h0);
  reg [(4'h8):(1'h0)] reg1241 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1239 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1238 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1237 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1236 = (1'h0);
  reg [(4'h9):(1'h0)] reg1232 = (1'h0);
  reg [(5'h18):(1'h0)] forvar1231 = (1'h0);
  reg [(4'h8):(1'h0)] forvar1230 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1226 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1220 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1219 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1218 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1217 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1215 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1214 = (1'h0);
  reg [(2'h2):(1'h0)] reg119 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg118 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar117 = (1'h0);
  reg [(4'he):(1'h0)] reg115 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg114 = (1'h0);
  reg [(4'he):(1'h0)] reg113 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg112 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg107 = (1'h0);
  reg [(4'hc):(1'h0)] forvar106 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar103 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg102 = (1'h0);
  reg [(4'h8):(1'h0)] reg98 = (1'h0);
  reg [(2'h2):(1'h0)] forvar96 = (1'h0);
  reg [(5'h18):(1'h0)] reg94 = (1'h0);
  reg [(3'h6):(1'h0)] reg90 = (1'h0);
  reg [(4'h9):(1'h0)] reg88 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg86 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar85 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg84 = (1'h0);
  reg [(3'h6):(1'h0)] reg80 = (1'h0);
  reg [(3'h6):(1'h0)] forvar79 = (1'h0);
  reg [(4'he):(1'h0)] reg77 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg76 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg73 = (1'h0);
  reg [(3'h5):(1'h0)] reg71 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar68 = (1'h0);
  reg [(4'h8):(1'h0)] reg66 = (1'h0);
  reg [(4'hc):(1'h0)] reg65 = (1'h0);
  reg [(4'hb):(1'h0)] reg64 = (1'h0);
  reg [(5'h14):(1'h0)] reg62 = (1'h0);
  reg [(2'h3):(1'h0)] forvar61 = (1'h0);
  reg [(5'h17):(1'h0)] reg60 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg59 = (1'h0);
  reg [(4'he):(1'h0)] reg58 = (1'h0);
  reg [(5'h17):(1'h0)] reg56 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg54 = (1'h0);
  reg [(5'h16):(1'h0)] reg53 = (1'h0);
  reg [(5'h17):(1'h0)] reg52 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg51 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg50 = (1'h0);
  reg [(4'hc):(1'h0)] reg48 = (1'h0);
  reg [(3'h4):(1'h0)] forvar47 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar46 = (1'h0);
  reg [(5'h11):(1'h0)] forvar39 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg38 = (1'h0);
  reg [(5'h15):(1'h0)] forvar36 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg35 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg28 = (1'h0);
  reg [(4'hc):(1'h0)] reg23 = (1'h0);
  reg [(5'h12):(1'h0)] reg20 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg33 = (1'h0);
  reg [(5'h13):(1'h0)] reg32 = (1'h0);
  reg [(5'h13):(1'h0)] reg30 = (1'h0);
  reg [(4'h8):(1'h0)] reg29 = (1'h0);
  reg [(4'hb):(1'h0)] forvar28 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg25 = (1'h0);
  reg [(4'hd):(1'h0)] reg24 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar23 = (1'h0);
  reg [(5'h15):(1'h0)] forvar20 = (1'h0);
  reg [(5'h14):(1'h0)] reg19 = (1'h0);
  reg [(5'h18):(1'h0)] reg18 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg12 = (1'h0);
  reg [(5'h14):(1'h0)] forvar10 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg9 = (1'h0);
  reg signed [(3'h7):(1'h0)] forvar8 = (1'h0);
  reg [(4'hc):(1'h0)] reg7 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar6 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg5 = (1'h0);
  assign y = {wire1389,
                 wire1388,
                 wire1342,
                 wire1336,
                 wire1335,
                 wire1291,
                 wire1290,
                 wire1261,
                 wire1260,
                 wire1211,
                 wire120,
                 wire4,
                 reg1392,
                 reg1387,
                 reg1384,
                 reg1382,
                 reg1379,
                 reg1378,
                 reg1376,
                 reg1375,
                 reg1374,
                 reg1372,
                 reg1370,
                 reg1368,
                 reg1365,
                 reg1356,
                 reg1355,
                 reg1354,
                 reg1351,
                 reg1350,
                 reg1348,
                 reg1347,
                 reg1344,
                 reg1341,
                 reg1337,
                 reg1334,
                 reg1332,
                 reg1331,
                 reg1330,
                 reg1327,
                 reg1323,
                 reg1321,
                 reg1320,
                 reg1314,
                 reg1311,
                 reg1307,
                 reg1306,
                 reg1305,
                 reg1303,
                 reg1300,
                 reg1296,
                 reg1295,
                 reg1292,
                 reg1286,
                 reg1281,
                 reg1278,
                 reg1277,
                 reg1276,
                 reg1274,
                 reg1271,
                 reg1269,
                 reg1267,
                 reg1266,
                 reg1263,
                 reg1259,
                 reg1255,
                 reg1254,
                 reg1246,
                 reg1245,
                 reg1242,
                 reg1240,
                 reg1235,
                 reg1234,
                 reg1233,
                 reg1229,
                 reg1228,
                 reg1227,
                 reg1225,
                 reg1224,
                 reg1223,
                 reg1222,
                 reg1221,
                 reg1216,
                 reg1213,
                 reg116,
                 reg111,
                 reg110,
                 reg109,
                 reg108,
                 reg105,
                 reg104,
                 reg101,
                 reg100,
                 reg99,
                 reg97,
                 reg95,
                 reg93,
                 reg92,
                 reg85,
                 reg91,
                 reg89,
                 reg87,
                 reg83,
                 reg82,
                 reg81,
                 reg78,
                 reg75,
                 reg74,
                 reg72,
                 reg70,
                 reg69,
                 reg67,
                 reg63,
                 reg57,
                 reg55,
                 reg49,
                 reg45,
                 reg44,
                 reg43,
                 reg42,
                 reg41,
                 reg40,
                 reg37,
                 reg34,
                 reg31,
                 reg27,
                 reg26,
                 reg22,
                 reg21,
                 reg17,
                 reg16,
                 reg15,
                 reg14,
                 reg13,
                 reg11,
                 reg1391,
                 reg1390,
                 reg1386,
                 forvar1385,
                 forvar1373,
                 forvar1368,
                 reg1383,
                 reg1381,
                 reg1380,
                 reg1377,
                 reg1373,
                 reg1371,
                 reg1369,
                 reg1367,
                 reg1366,
                 reg1364,
                 reg1363,
                 forvar1362,
                 reg1361,
                 forvar1360,
                 reg1359,
                 reg1358,
                 reg1357,
                 forvar1354,
                 reg1352,
                 reg1353,
                 forvar1352,
                 forvar1349,
                 reg1343,
                 reg1346,
                 reg1345,
                 forvar1343,
                 reg1340,
                 reg1339,
                 reg1338,
                 reg1333,
                 reg1329,
                 reg1328,
                 reg1326,
                 reg1325,
                 reg1324,
                 reg1322,
                 forvar1319,
                 reg1318,
                 reg1317,
                 reg1316,
                 reg1315,
                 forvar1313,
                 reg1312,
                 reg1310,
                 reg1309,
                 forvar1308,
                 reg1304,
                 reg1302,
                 reg1301,
                 reg1299,
                 reg1298,
                 reg1293,
                 forvar1292,
                 reg1297,
                 reg1294,
                 forvar1293,
                 reg1289,
                 reg1288,
                 reg1287,
                 reg1285,
                 forvar1284,
                 reg1283,
                 forvar1282,
                 reg1280,
                 reg1279,
                 forvar1275,
                 reg1273,
                 reg1272,
                 forvar1270,
                 forvar1268,
                 reg1265,
                 reg1264,
                 forvar1262,
                 reg1258,
                 reg1257,
                 reg1256,
                 forvar1253,
                 reg1252,
                 reg1251,
                 forvar1250,
                 forvar1249,
                 reg1248,
                 reg1247,
                 reg1244,
                 reg1243,
                 reg1241,
                 reg1239,
                 reg1238,
                 reg1237,
                 forvar1236,
                 reg1232,
                 forvar1231,
                 forvar1230,
                 reg1226,
                 reg1220,
                 reg1219,
                 reg1218,
                 reg1217,
                 forvar1215,
                 forvar1214,
                 reg119,
                 reg118,
                 forvar117,
                 reg115,
                 reg114,
                 reg113,
                 reg112,
                 reg107,
                 forvar106,
                 forvar103,
                 reg102,
                 reg98,
                 forvar96,
                 reg94,
                 reg90,
                 reg88,
                 reg86,
                 forvar85,
                 reg84,
                 reg80,
                 forvar79,
                 reg77,
                 reg76,
                 reg73,
                 reg71,
                 forvar68,
                 reg66,
                 reg65,
                 reg64,
                 reg62,
                 forvar61,
                 reg60,
                 reg59,
                 reg58,
                 reg56,
                 reg54,
                 reg53,
                 reg52,
                 reg51,
                 reg50,
                 reg48,
                 forvar47,
                 forvar46,
                 forvar39,
                 reg38,
                 forvar36,
                 reg35,
                 reg28,
                 reg23,
                 reg20,
                 reg33,
                 reg32,
                 reg30,
                 reg29,
                 forvar28,
                 reg25,
                 reg24,
                 forvar23,
                 forvar20,
                 reg19,
                 reg18,
                 reg12,
                 forvar10,
                 reg9,
                 forvar8,
                 reg7,
                 forvar6,
                 reg5,
                 (1'h0)};
  assign wire4 = (|(({(&wire1)} > wire3) ?
                     wire0[(4'hd):(4'h9)] : $unsigned($unsigned((-wire1)))));
  always
    @(posedge clk) begin
      reg5 = wire1;
      for (forvar6 = (1'h0); (forvar6 < (1'h0)); forvar6 = (forvar6 + (1'h1)))
        begin
          reg7 = (wire0[(4'h9):(2'h2)] ?
              forvar6[(3'h5):(1'h0)] : wire0[(5'h10):(3'h6)]);
          for (forvar8 = (1'h0); (forvar8 < (3'h4)); forvar8 = (forvar8 + (1'h1)))
            begin
              reg9 = $unsigned((~$unsigned((wire4 << (^~wire0)))));
            end
          for (forvar10 = (1'h0); (forvar10 < (3'h4)); forvar10 = (forvar10 + (1'h1)))
            begin
              reg11 <= ($unsigned(wire4[(2'h3):(1'h1)]) && wire0);
              reg12 = $signed($signed($signed((wire1 ?
                  $unsigned(wire4) : (!forvar8)))));
              reg13 <= forvar8;
              reg14 <= ((+$signed($unsigned(wire2))) ?
                  $unsigned(forvar8[(3'h4):(3'h4)]) : reg11[(4'h8):(1'h1)]);
            end
          reg15 <= (~&$signed(reg5[(2'h2):(1'h0)]));
          if ((8'hb8))
            begin
              reg16 <= (($signed((~|reg9)) && (!$signed($signed(reg7)))) || {$signed($signed(reg11[(3'h7):(2'h2)])),
                  $signed(wire2)});
              reg17 <= ($signed($unsigned((!reg7[(4'h9):(3'h5)]))) < $signed(({(reg11 ?
                      wire1 : reg14),
                  {wire1, reg14}} >>> $signed((+forvar6)))));
              reg18 = (|$signed(((~&reg13[(4'hb):(2'h2)]) ? wire0 : reg7)));
            end
          else
            begin
              reg16 <= $signed((~|(~&((&reg16) ?
                  (|reg13) : $unsigned(reg13)))));
              reg17 <= wire0;
              reg18 = ({{((reg11 ? wire1 : (8'hb5)) >= (~^reg11)),
                          (forvar8[(3'h4):(2'h2)] ?
                              $signed(reg14) : (~|reg18))},
                      $signed($signed($unsigned(wire1)))} ?
                  reg14 : wire2[(1'h0):(1'h0)]);
            end
        end
      reg19 = (wire3[(4'h8):(4'h8)] ? wire3 : $unsigned(wire2));
    end
  always
    @(posedge clk) begin
      if ($unsigned($unsigned(((~|{reg13, reg17}) ?
          reg15 : reg16[(3'h7):(1'h1)]))))
        begin
          for (forvar20 = (1'h0); (forvar20 < (2'h2)); forvar20 = (forvar20 + (1'h1)))
            begin
              reg21 <= ((($signed(wire3) ?
                      ($signed((8'hab)) < (8'ha7)) : reg17[(2'h2):(2'h2)]) ?
                  wire3 : $signed($unsigned($signed((8'ha1))))) | (^~{$signed(reg17[(1'h1):(1'h0)])}));
              reg22 <= ({(reg16[(1'h0):(1'h0)] ?
                          ((reg11 != (8'hb2)) ~^ reg17[(2'h2):(1'h0)]) : forvar20),
                      (~^reg15[(4'hb):(1'h0)])} ?
                  (8'hbb) : $unsigned($unsigned($signed($unsigned(reg14)))));
            end
          for (forvar23 = (1'h0); (forvar23 < (2'h3)); forvar23 = (forvar23 + (1'h1)))
            begin
              reg24 = $signed(reg11);
              reg25 = ({(+reg16[(3'h6):(2'h2)]), forvar23[(4'hb):(4'h8)]} ?
                  reg16[(2'h3):(1'h1)] : forvar20);
              reg26 <= ((|{$signed((7'h47))}) || $signed({$unsigned(reg17),
                  ($signed(wire2) ? $signed((8'ha1)) : {reg11})}));
              reg27 <= {(({$unsigned(reg16), (reg11 && forvar20)} != (reg15 ?
                          reg17 : wire3[(4'he):(4'hc)])) ?
                      forvar23 : $unsigned(((wire2 ? (8'hb5) : (8'ha9)) ?
                          reg22 : reg15[(1'h0):(1'h0)]))),
                  ($signed($signed($signed(wire2))) ?
                      (reg21[(2'h3):(1'h0)] ?
                          (reg26[(5'h15):(5'h13)] > reg11) : ((|reg17) ?
                              $unsigned(forvar23) : (forvar20 && wire2))) : ((~&{reg11,
                              reg14}) ?
                          ({wire3, reg15} | $signed(reg25)) : reg26))};
            end
          for (forvar28 = (1'h0); (forvar28 < (1'h0)); forvar28 = (forvar28 + (1'h1)))
            begin
              reg29 = reg17;
              reg30 = (-reg14[(4'hd):(2'h3)]);
              reg31 <= wire0;
              reg32 = reg26;
              reg33 = wire1;
            end
        end
      else
        begin
          reg20 = ((((!(reg27 ? (8'hb4) : reg33)) ?
                  (reg25 <<< $unsigned(reg33)) : (^$signed(reg32))) ?
              (~$signed({reg13, reg25})) : forvar20[(3'h6):(1'h1)]) <<< (reg17 ?
              wire4[(4'hb):(4'hb)] : reg26[(3'h6):(3'h6)]));
          if (($unsigned((reg30[(4'hb):(3'h6)] <<< ({(8'ha9)} && ((8'ha0) || reg25)))) * $unsigned(reg13)))
            begin
              reg23 = wire3;
            end
          else
            begin
              reg23 = ($unsigned(reg20) < (~^(~^$signed((reg25 ?
                  (8'hb4) : reg23)))));
              reg26 <= $unsigned((!($signed({reg17, reg32}) ^~ ((^~reg33) ?
                  $signed((8'hb9)) : $signed(wire2)))));
              reg27 <= ((reg33 ?
                      (($signed((7'h45)) ^~ $unsigned(reg22)) ?
                          ((reg15 ? reg20 : reg24) ?
                              (reg21 < reg15) : (~&forvar20)) : $signed((reg16 <<< (8'hbc)))) : (reg33 != (~^reg25))) ?
                  (($signed((reg29 ? reg14 : reg13)) >> ((reg14 ?
                              reg26 : wire2) ?
                          (reg16 != wire2) : (reg11 << reg25))) ?
                      ({((8'ha0) >> reg26)} | $signed((&forvar28))) : $signed(forvar28[(4'h9):(1'h0)])) : reg14);
              reg28 = reg32[(4'hb):(3'h5)];
              reg31 <= reg17;
            end
          reg34 <= $unsigned(reg17);
          reg35 = $unsigned({$unsigned(reg26[(4'ha):(3'h7)]),
              $signed(wire1[(2'h3):(2'h3)])});
        end
      for (forvar36 = (1'h0); (forvar36 < (2'h2)); forvar36 = (forvar36 + (1'h1)))
        begin
          reg37 <= (((8'ha7) ? (^~reg29[(3'h7):(3'h5)]) : reg21) ^ forvar23);
          reg38 = {$unsigned($unsigned((reg34 ?
                  {forvar23, (8'h9c)} : (reg33 ? forvar20 : reg27)))),
              $unsigned((-(8'ha7)))};
          for (forvar39 = (1'h0); (forvar39 < (2'h2)); forvar39 = (forvar39 + (1'h1)))
            begin
              reg40 <= {(~^$unsigned(reg26[(5'h15):(5'h15)])),
                  (forvar20 ?
                      (reg26[(1'h0):(1'h0)] >= ((8'ha4) ~^ $signed(reg32))) : $signed($signed(((8'ha5) ?
                          reg28 : reg17))))};
              reg41 <= $unsigned((8'hbb));
              reg42 <= (($unsigned((~^((7'h48) <<< reg17))) != (forvar20 ?
                  forvar28[(3'h6):(1'h1)] : ({reg38,
                      forvar39} && (~^wire2)))) | ((reg24 ?
                  $unsigned((~^reg33)) : {(-reg37)}) >>> ((8'hb1) ?
                  (~$signed(reg35)) : (reg23 ? reg22 : reg20[(3'h6):(1'h0)]))));
              reg43 <= (~^$signed(reg41));
            end
          reg44 <= (~^$unsigned({reg26}));
        end
      reg45 <= (wire4 ? reg31[(3'h6):(3'h5)] : forvar36);
    end
  always
    @(posedge clk) begin
      for (forvar46 = (1'h0); (forvar46 < (2'h3)); forvar46 = (forvar46 + (1'h1)))
        begin
          for (forvar47 = (1'h0); (forvar47 < (1'h0)); forvar47 = (forvar47 + (1'h1)))
            begin
              reg48 = reg45;
            end
          reg49 <= $signed((($unsigned((!reg11)) ? reg41 : reg26) ?
              reg17[(1'h0):(1'h0)] : $signed(wire2[(3'h7):(2'h3)])));
          reg50 = reg41[(5'h11):(5'h10)];
          if ((~{$unsigned((|reg15)), reg22}))
            begin
              reg51 = $unsigned($signed((((-reg41) && (reg43 - wire0)) ?
                  $signed($unsigned(reg16)) : $unsigned((forvar46 >> reg15)))));
              reg52 = $signed(reg50);
            end
          else
            begin
              reg51 = $signed(reg16);
              reg52 = $unsigned((~|$unsigned(reg52[(4'hb):(3'h6)])));
              reg53 = (8'hb7);
              reg54 = {reg27,
                  (((^$unsigned(reg50)) ?
                          reg43 : (reg22[(1'h1):(1'h0)] * $signed(reg51))) ?
                      (&$unsigned($signed(reg26))) : (reg22 ?
                          (|reg45) : reg31[(4'hd):(2'h2)]))};
              reg55 <= reg54;
            end
          if (reg37)
            begin
              reg56 = reg26;
              reg57 <= (~|$unsigned({(~|$unsigned(wire2)),
                  (^$unsigned(reg40))}));
              reg58 = {{(reg31 ? $signed((+reg56)) : reg43),
                      $unsigned($signed((8'ha7)))}};
              reg59 = (!$signed((forvar47[(1'h1):(1'h1)] ?
                  $signed((|reg14)) : $unsigned(((8'h9f) <= wire1)))));
              reg60 = {reg52[(3'h7):(1'h0)]};
            end
          else
            begin
              reg57 <= $signed($unsigned(($unsigned(reg42[(3'h4):(2'h3)]) || ((wire0 <<< reg42) >> $unsigned(reg15)))));
            end
        end
      for (forvar61 = (1'h0); (forvar61 < (1'h0)); forvar61 = (forvar61 + (1'h1)))
        begin
          if (({wire3, $unsigned(reg49)} ?
              $unsigned(reg49[(3'h5):(1'h0)]) : reg43[(1'h0):(1'h0)]))
            begin
              reg62 = {reg11[(3'h7):(3'h4)],
                  (reg60 ^ $unsigned($unsigned($unsigned(reg15))))};
            end
          else
            begin
              reg63 <= (reg53 || (~(~|forvar61)));
              reg64 = reg26;
              reg65 = reg57;
              reg66 = (!$signed(wire4));
              reg67 <= reg50;
            end
          for (forvar68 = (1'h0); (forvar68 < (1'h1)); forvar68 = (forvar68 + (1'h1)))
            begin
              reg69 <= (&(8'hb2));
              reg70 <= reg17;
              reg71 = reg17[(2'h2):(1'h1)];
              reg72 <= $unsigned((forvar68 ?
                  reg50[(2'h3):(2'h3)] : (reg49[(1'h0):(1'h0)] && ((reg11 ?
                      (8'hb0) : (8'hbc)) + {reg22, wire2}))));
            end
          reg73 = (+((~(reg41 ?
              (reg50 >> reg22) : $signed(reg69))) * ({reg70} >>> reg62[(4'hc):(1'h0)])));
          if (((~&$signed($unsigned((reg15 ? reg34 : reg11)))) ?
              reg65[(3'h5):(1'h0)] : reg59))
            begin
              reg74 <= (~^((((~^reg27) ? $unsigned(reg17) : reg51) ?
                  (~^$unsigned(reg52)) : {reg51[(2'h2):(2'h2)],
                      reg43[(4'h9):(2'h2)]}) <= (reg17[(1'h0):(1'h0)] ?
                  $signed((8'h9d)) : forvar68[(4'hf):(4'he)])));
              reg75 <= $unsigned(reg50);
            end
          else
            begin
              reg74 <= ({($unsigned(reg42) ?
                          ($unsigned(reg62) ?
                              wire1[(4'hf):(4'hf)] : ((8'ha4) >>> reg52)) : ($signed((8'hbe)) ?
                              $signed(reg67) : ((7'h45) ? (8'hb0) : wire0)))} ?
                  ({reg58, $unsigned({wire0, wire0})} ?
                      $unsigned(reg58[(1'h0):(1'h0)]) : (reg75 ~^ (-$signed(reg72)))) : $signed((8'had)));
              reg76 = reg40[(3'h6):(2'h2)];
              reg77 = reg26[(5'h12):(4'h8)];
              reg78 <= (-$unsigned($signed(reg50)));
            end
          for (forvar79 = (1'h0); (forvar79 < (2'h2)); forvar79 = (forvar79 + (1'h1)))
            begin
              reg80 = ($unsigned(reg45) - $unsigned($signed((reg15[(4'ha):(3'h6)] >> $signed(reg71)))));
              reg81 <= (8'hb2);
              reg82 <= (&$unsigned({(reg73 ?
                      (reg70 ? reg64 : reg81) : (reg60 | reg59)),
                  reg41}));
            end
        end
      reg83 <= reg67[(3'h4):(3'h4)];
      reg84 = ($signed(reg62) ? reg82 : reg64);
    end
  always
    @(posedge clk) begin
      if ((-{$unsigned(reg69), reg70[(1'h0):(1'h0)]}))
        begin
          for (forvar85 = (1'h0); (forvar85 < (1'h1)); forvar85 = (forvar85 + (1'h1)))
            begin
              reg86 = $unsigned($signed(((((8'haf) ?
                      reg55 : reg42) - $unsigned((8'ha8))) ?
                  reg78[(3'h7):(3'h5)] : ((reg45 - reg72) > $signed((8'hb1))))));
              reg87 <= (~&reg31[(3'h7):(1'h0)]);
              reg88 = $signed((8'haf));
            end
          reg89 <= ($unsigned($signed($signed((reg43 ?
              reg37 : reg43)))) <<< ((^((~reg22) ?
                  (reg22 ? reg34 : (8'haa)) : $signed(reg42))) ?
              {((8'hae) << (reg67 ? reg88 : reg37))} : (((reg44 || reg31) ?
                  $unsigned(reg37) : wire2[(4'hc):(2'h2)]) >>> (reg70 ?
                  (~reg57) : reg11[(4'he):(4'h8)]))));
          reg90 = (-((reg34 ~^ (^~(reg14 ? reg41 : reg42))) <= reg45));
          reg91 <= (8'hb8);
        end
      else
        begin
          reg85 <= (~$unsigned(reg40[(5'h10):(4'hd)]));
          if (reg42)
            begin
              reg87 <= {$unsigned((~(reg11[(5'h10):(4'hd)] >> reg72)))};
              reg88 = (reg87 ?
                  (($unsigned($signed(reg70)) || (~^(reg42 ?
                      (8'haa) : reg70))) ^ ((&(+reg41)) | reg31)) : {(|((reg42 == (8'hab)) ?
                          $unsigned(reg74) : {reg42, reg16})),
                      ((reg26[(3'h7):(2'h2)] != $signed(reg44)) >>> ((~|reg85) ^~ (^reg14)))});
              reg89 <= (8'hbb);
              reg91 <= (($signed(((reg31 * reg75) ?
                      (~^reg75) : $unsigned(reg72))) ?
                  $signed({wire4,
                      reg72}) : reg14) >>> ($signed((+reg27)) | $unsigned($unsigned(reg88[(2'h3):(1'h1)]))));
              reg92 <= reg13;
            end
          else
            begin
              reg87 <= (reg75 ?
                  $signed($signed($unsigned(reg81))) : $unsigned((-$unsigned($signed(reg82)))));
              reg89 <= reg63[(4'hb):(3'h4)];
            end
          if (reg43[(3'h5):(2'h2)])
            begin
              reg93 <= reg31;
            end
          else
            begin
              reg93 <= ((((~|(^reg17)) ?
                  wire0[(4'h9):(3'h4)] : reg43) != (~&$signed((reg82 >> reg82)))) < reg45);
              reg94 = $signed((reg69[(5'h13):(4'hf)] || reg69[(1'h0):(1'h0)]));
              reg95 <= (+({reg63[(3'h4):(1'h1)]} ?
                  (8'haf) : (reg75 ? (^$unsigned(reg21)) : (!(~&reg63)))));
            end
          for (forvar96 = (1'h0); (forvar96 < (3'h4)); forvar96 = (forvar96 + (1'h1)))
            begin
              reg97 <= wire1[(1'h0):(1'h0)];
              reg98 = $signed(reg97[(3'h4):(2'h3)]);
              reg99 <= $unsigned((+$signed((reg13[(1'h1):(1'h0)] >>> {wire0}))));
            end
          reg100 <= (($unsigned($unsigned((-(8'ha3)))) & ((reg81 | (8'had)) ~^ $signed($unsigned(wire4)))) >= ($signed(($unsigned((8'had)) ?
                  $signed(reg42) : (&reg89))) ?
              ($signed({reg45}) ?
                  reg78[(4'h8):(1'h1)] : $signed((8'hb8))) : reg15[(5'h15):(5'h15)]));
        end
      reg101 <= $unsigned($signed(reg15[(5'h12):(3'h5)]));
      reg102 = ({($signed((reg34 ^ forvar96)) ? reg57 : reg41)} ?
          $signed($unsigned($unsigned((reg100 ? reg72 : reg43)))) : reg11);
      for (forvar103 = (1'h0); (forvar103 < (2'h2)); forvar103 = (forvar103 + (1'h1)))
        begin
          reg104 <= (reg69 << reg55[(4'ha):(1'h0)]);
          reg105 <= (($signed((~&$signed(wire2))) ?
              (~reg75[(4'ha):(3'h7)]) : reg104[(4'h9):(3'h4)]) >= {((forvar85[(4'h8):(1'h0)] ?
                  (reg15 - reg89) : ((8'ha2) <= (8'haa))) <= (&$signed(reg97)))});
          for (forvar106 = (1'h0); (forvar106 < (1'h0)); forvar106 = (forvar106 + (1'h1)))
            begin
              reg107 = $signed(((reg70[(2'h3):(1'h0)] ?
                      $signed((wire2 != forvar96)) : $signed($unsigned(reg78))) ?
                  wire3 : (~|((|reg15) << (8'hbb)))));
              reg108 <= (((|wire0) ?
                      ($unsigned(reg26[(5'h13):(3'h6)]) ^ {$unsigned((7'h45))}) : ($unsigned((~|reg26)) ?
                          {(reg11 - reg72),
                              (reg13 || reg78)} : (reg97 >>> (+reg107)))) ?
                  (~^$signed($signed((~&(8'hac))))) : $unsigned(reg72[(3'h7):(3'h7)]));
              reg109 <= $unsigned($signed(((reg55 ?
                  reg74 : (reg21 <= reg88)) ~^ $signed((reg67 ^ wire4)))));
              reg110 <= (({(-$unsigned(reg69))} ?
                  ($unsigned(reg49[(4'he):(2'h3)]) ?
                      $signed(reg22[(2'h3):(1'h0)]) : $unsigned($signed(reg95))) : reg63[(4'hb):(2'h3)]) < {forvar85[(1'h0):(1'h0)]});
              reg111 <= $signed({(~^(^~{reg72, reg101}))});
            end
          if ({{(~((~reg13) ? {reg108, reg102} : (wire1 ? reg98 : (7'h47))))}})
            begin
              reg112 = wire3;
              reg113 = $signed(reg74);
              reg114 = ((reg78[(2'h2):(1'h1)] | ($signed($signed((8'hbe))) ?
                      reg97 : ((7'h4a) ? reg22[(1'h1):(1'h0)] : reg11))) ?
                  (|(8'hb0)) : (~^(~{{reg86}, (&reg86)})));
              reg115 = (($signed((8'hb0)) ?
                      reg49[(3'h4):(1'h0)] : $unsigned(reg70[(2'h2):(2'h2)])) ?
                  reg112 : (~wire2[(5'h14):(1'h1)]));
              reg116 <= $signed((&{$signed((~reg74)), $unsigned((-wire3))}));
            end
          else
            begin
              reg112 = $unsigned({(~|((~^reg22) ?
                      reg98[(3'h7):(2'h3)] : (reg82 == reg31))),
                  (+$signed($unsigned(reg67)))});
              reg116 <= $unsigned($unsigned({(reg87 > reg81[(1'h1):(1'h0)])}));
            end
          for (forvar117 = (1'h0); (forvar117 < (2'h2)); forvar117 = (forvar117 + (1'h1)))
            begin
              reg118 = forvar106[(4'hb):(1'h0)];
              reg119 = $unsigned($unsigned($signed((|reg67))));
            end
        end
    end
  assign wire120 = $unsigned($unsigned((^~(7'h47))));
  module121 #() modinst1212 (.wire124(reg82), .y(wire1211), .wire125(reg101), .wire122(reg16), .wire123(reg72), .clk(clk));
  always
    @(posedge clk) begin
      reg1213 <= $unsigned($unsigned(reg37[(2'h2):(1'h0)]));
      for (forvar1214 = (1'h0); (forvar1214 < (2'h3)); forvar1214 = (forvar1214 + (1'h1)))
        begin
          for (forvar1215 = (1'h0); (forvar1215 < (2'h3)); forvar1215 = (forvar1215 + (1'h1)))
            begin
              reg1216 <= (reg14[(4'he):(4'hb)] < reg11);
              reg1217 = $signed($signed(reg87));
              reg1218 = reg1216[(4'h8):(2'h2)];
              reg1219 = ((((reg21 >>> (reg49 ? reg85 : reg104)) ?
                      ($unsigned(reg82) ?
                          $unsigned(reg70) : (reg99 ?
                              reg21 : reg17)) : reg87[(5'h10):(4'hc)]) ?
                  $signed(reg105[(4'ha):(3'h4)]) : $signed(reg22[(2'h2):(1'h0)])) - reg43[(4'ha):(3'h5)]);
              reg1220 = reg1217[(1'h0):(1'h0)];
            end
          if (reg14[(3'h4):(2'h3)])
            begin
              reg1221 <= reg26[(4'he):(4'he)];
              reg1222 <= reg97;
              reg1223 <= (~^(~&$unsigned(((|reg45) == reg57[(2'h3):(1'h1)]))));
              reg1224 <= $unsigned($signed(reg37[(2'h3):(2'h3)]));
              reg1225 <= (({$signed(reg49), $signed((reg16 ? reg31 : reg87))} ?
                      $signed(reg31) : $signed(((reg63 >>> reg75) && (reg100 * reg67)))) ?
                  $signed(({$signed(reg63)} ?
                      reg1213[(2'h2):(1'h0)] : reg11[(5'h17):(3'h7)])) : (|$unsigned(($unsigned(reg92) ?
                      reg40[(4'hb):(4'h8)] : (reg83 << reg1219)))));
            end
          else
            begin
              reg1221 <= $signed(($signed(reg1221[(3'h6):(2'h2)]) != reg45));
              reg1226 = reg75;
              reg1227 <= $signed(reg91[(4'hd):(3'h4)]);
            end
        end
      reg1228 <= {$unsigned(((|(reg99 && reg1220)) || ($signed(reg116) ^ $unsigned(wire4)))),
          {wire4[(2'h3):(2'h2)],
              (reg87 ?
                  $unsigned(reg1221) : {(reg1222 << reg111),
                      (reg11 <<< reg1220)})}};
      reg1229 <= (reg31 ?
          (~|$unsigned((reg63[(4'ha):(3'h4)] && (reg83 ?
              reg104 : reg44)))) : $signed($signed(reg67[(4'h8):(3'h7)])));
      for (forvar1230 = (1'h0); (forvar1230 < (1'h0)); forvar1230 = (forvar1230 + (1'h1)))
        begin
          for (forvar1231 = (1'h0); (forvar1231 < (3'h4)); forvar1231 = (forvar1231 + (1'h1)))
            begin
              reg1232 = reg111[(1'h1):(1'h0)];
              reg1233 <= (8'hb3);
              reg1234 <= $signed(wire2[(4'hb):(3'h4)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg1235 <= reg1223[(5'h11):(1'h0)];
      for (forvar1236 = (1'h0); (forvar1236 < (2'h2)); forvar1236 = (forvar1236 + (1'h1)))
        begin
          reg1237 = $signed($signed(wire4));
          if (({(-reg67[(1'h0):(1'h0)])} && (&(~&{$signed(reg109)}))))
            begin
              reg1238 = (~&$signed(((+{reg1237}) <<< reg42[(2'h2):(2'h2)])));
              reg1239 = ((!reg26) && $signed($unsigned(((reg104 ?
                  reg87 : reg1213) ^ ((8'hae) ? reg105 : reg1229)))));
              reg1240 <= ((!($unsigned($unsigned(reg1237)) > ((reg69 ^~ (8'hb4)) ?
                      (wire3 << reg43) : (reg75 ? wire3 : reg21)))) ?
                  $signed($unsigned((+(reg1228 | wire1)))) : reg69[(5'h12):(4'hd)]);
              reg1241 = ($signed(((reg92[(4'h9):(3'h6)] ?
                          (reg1238 < reg43) : reg116) ?
                      (7'h45) : (~&$unsigned(reg14)))) ?
                  (reg1228 ?
                      (reg27[(4'hb):(3'h6)] ~^ reg1233[(3'h4):(2'h2)]) : (-$signed((reg95 >= (8'hb3))))) : $signed(($unsigned(reg13[(3'h7):(3'h4)]) >= (wire1[(4'hf):(4'h8)] ?
                      $signed(reg17) : reg44[(5'h14):(5'h12)]))));
            end
          else
            begin
              reg1240 <= (reg69 > reg44);
            end
          reg1242 <= reg111;
          if ($signed(wire4))
            begin
              reg1243 = (((~^($signed(wire0) ~^ (reg74 ?
                  reg108 : reg40))) * reg43[(3'h6):(3'h5)]) ~^ (-reg1225));
              reg1244 = wire3[(3'h5):(3'h5)];
            end
          else
            begin
              reg1245 <= reg1243;
              reg1246 <= $unsigned(reg21);
              reg1247 = ((^(~&$signed({reg37, wire4}))) << ((7'h43) >>> reg49));
              reg1248 = $signed((&{$unsigned($signed(reg110)), reg100}));
            end
        end
      for (forvar1249 = (1'h0); (forvar1249 < (1'h1)); forvar1249 = (forvar1249 + (1'h1)))
        begin
          for (forvar1250 = (1'h0); (forvar1250 < (1'h0)); forvar1250 = (forvar1250 + (1'h1)))
            begin
              reg1251 = (~&$signed({reg91}));
            end
          reg1252 = reg1224;
          for (forvar1253 = (1'h0); (forvar1253 < (3'h4)); forvar1253 = (forvar1253 + (1'h1)))
            begin
              reg1254 <= {($signed($signed($unsigned(reg67))) ~^ ((reg1235[(1'h0):(1'h0)] ?
                          (reg1229 ? (8'hbc) : reg1216) : (reg1225 ?
                              (8'hb3) : reg101)) ?
                      $signed((reg1233 ? reg11 : reg99)) : reg1240)),
                  (!(((|(8'h9e)) ?
                      $signed((8'ha6)) : (reg99 & reg1221)) > $unsigned((reg81 ?
                      reg92 : reg1252))))};
              reg1255 <= (($signed(reg41[(3'h5):(1'h0)]) ?
                  ((~(~reg1235)) ?
                      ($signed(reg1233) ?
                          (8'ha7) : ((8'hb8) & reg99)) : ((reg78 ~^ reg1254) << (^~reg22))) : {reg1243}) > reg42);
              reg1256 = $unsigned($signed(reg22));
            end
          reg1257 = (~|$unsigned((-($signed(reg15) ?
              reg93 : $signed(forvar1236)))));
        end
      reg1258 = $signed((|($unsigned(reg27) ?
          (^~(forvar1253 ? reg13 : reg108)) : reg1251[(5'h12):(5'h11)])));
      reg1259 <= reg104[(3'h6):(3'h4)];
    end
  assign wire1260 = $signed(reg105);
  assign wire1261 = reg43[(4'hb):(3'h4)];
  always
    @(posedge clk) begin
      for (forvar1262 = (1'h0); (forvar1262 < (2'h3)); forvar1262 = (forvar1262 + (1'h1)))
        begin
          reg1263 <= (&(^{(reg109 ? $signed(reg1240) : reg22),
              $unsigned((reg21 ? reg69 : reg108))}));
          if (reg82[(1'h1):(1'h0)])
            begin
              reg1264 = $signed({((reg1227[(3'h6):(1'h0)] == reg17[(2'h3):(2'h2)]) ?
                      (7'h47) : {(reg91 ? (8'ha2) : (8'ha9))}),
                  wire1211});
              reg1265 = reg1224[(2'h2):(1'h0)];
            end
          else
            begin
              reg1266 <= $signed(((reg40 ?
                      {(reg91 ? reg1242 : reg1264)} : {(wire0 + (8'hae)),
                          (reg83 != reg105)}) ?
                  (^~$unsigned((reg70 >= (8'hb7)))) : (reg41 | (^~(+(8'ha2))))));
            end
          reg1267 <= ($signed({reg45[(2'h3):(2'h3)]}) ?
              (^(&reg15)) : $unsigned(($unsigned((~&reg1245)) ?
                  $unsigned(wire1260[(4'he):(4'ha)]) : ({reg1228} ?
                      reg95 : (+wire0)))));
        end
      for (forvar1268 = (1'h0); (forvar1268 < (3'h4)); forvar1268 = (forvar1268 + (1'h1)))
        begin
          reg1269 <= $unsigned((^~(reg97[(4'hc):(4'hb)] ?
              ((reg1245 ^ reg108) ?
                  (wire4 ? reg82 : reg1240) : ((8'hbc) ?
                      reg81 : wire2)) : (&$unsigned((7'h42))))));
          for (forvar1270 = (1'h0); (forvar1270 < (2'h2)); forvar1270 = (forvar1270 + (1'h1)))
            begin
              reg1271 <= ((~^{{$signed(reg1255), (reg109 == reg17)}}) ?
                  reg1221 : reg101);
              reg1272 = (((~($unsigned(reg91) ?
                      (reg13 ? reg1259 : reg55) : (^~reg67))) ?
                  forvar1268 : $signed(forvar1268[(2'h2):(1'h0)])) << reg1269);
              reg1273 = $unsigned(reg101);
            end
          reg1274 <= $unsigned(reg74[(5'h13):(4'h8)]);
          for (forvar1275 = (1'h0); (forvar1275 < (2'h3)); forvar1275 = (forvar1275 + (1'h1)))
            begin
              reg1276 <= (reg1266[(3'h7):(3'h6)] ?
                  {((~reg89) ?
                          {$unsigned(reg1255)} : $signed((reg1255 ?
                              reg16 : reg1234))),
                      $unsigned($signed(wire4[(2'h2):(1'h1)]))} : reg92[(4'h8):(1'h0)]);
              reg1277 <= {reg110, $unsigned(reg45[(1'h0):(1'h0)])};
              reg1278 <= wire3[(4'h8):(1'h1)];
              reg1279 = reg1255[(3'h5):(3'h5)];
              reg1280 = $signed(reg1278);
            end
          reg1281 <= (&$signed($signed($unsigned((reg83 >> reg1242)))));
        end
      for (forvar1282 = (1'h0); (forvar1282 < (3'h4)); forvar1282 = (forvar1282 + (1'h1)))
        begin
          reg1283 = ({reg1269,
              wire120[(1'h0):(1'h0)]} >> ((-$signed($unsigned(reg43))) & $unsigned($signed((~^reg95)))));
          for (forvar1284 = (1'h0); (forvar1284 < (1'h1)); forvar1284 = (forvar1284 + (1'h1)))
            begin
              reg1285 = forvar1262;
            end
          if ({$unsigned({(!(~&reg44)), $signed($signed(reg1265))})})
            begin
              reg1286 <= ($signed(reg21) ?
                  reg1246[(3'h5):(1'h0)] : $signed((|(~&(&(7'h41))))));
            end
          else
            begin
              reg1287 = reg1265[(3'h4):(2'h3)];
              reg1288 = (reg69[(4'ha):(2'h2)] ?
                  (reg14 ? (&reg63) : (8'ha2)) : ((|$unsigned(reg1278)) ?
                      reg72[(1'h0):(1'h0)] : reg108[(1'h0):(1'h0)]));
            end
          reg1289 = (^~(wire1[(1'h1):(1'h0)] <<< (reg31[(4'hc):(4'hb)] ?
              wire3[(4'hb):(3'h6)] : reg1283)));
        end
    end
  assign wire1290 = $unsigned(wire1260[(2'h3):(1'h0)]);
  assign wire1291 = reg21;
  always
    @(posedge clk) begin
      if (wire1)
        begin
          reg1292 <= (~|(|reg85));
          for (forvar1293 = (1'h0); (forvar1293 < (2'h3)); forvar1293 = (forvar1293 + (1'h1)))
            begin
              reg1294 = reg1213;
              reg1295 <= reg83[(1'h0):(1'h0)];
              reg1296 <= (reg34 << $signed(((~&(reg72 ?
                  reg1277 : reg1295)) ^ ($signed(reg14) == reg1281))));
              reg1297 = $signed(((((reg41 > (8'hb8)) >> $signed((7'h43))) <<< (reg99 << reg1228)) ^ reg87));
            end
        end
      else
        begin
          for (forvar1292 = (1'h0); (forvar1292 < (3'h4)); forvar1292 = (forvar1292 + (1'h1)))
            begin
              reg1293 = $signed($signed(wire1260));
              reg1295 <= (&(^~((7'h48) ?
                  {(~&reg1221)} : {$unsigned(reg1276)})));
            end
        end
      reg1298 = ($signed(($signed((reg1296 > reg1221)) & (reg78[(1'h0):(1'h0)] >> (|reg92)))) ?
          $unsigned(((~^reg1263[(1'h0):(1'h0)]) ?
              (~&$unsigned(reg1294)) : (|(reg1221 ^ reg1242)))) : reg22[(3'h4):(2'h3)]);
      if (reg27[(3'h6):(1'h0)])
        begin
          reg1299 = (reg55 ?
              (~&(^((reg1240 ? reg1228 : reg27) ?
                  reg63[(4'ha):(3'h7)] : $signed(reg1234)))) : $signed((~|((reg70 ?
                      reg1267 : forvar1292) ?
                  reg1221[(3'h6):(2'h2)] : reg85))));
          if (((($signed((&reg95)) ?
                      $signed({reg45, (7'h48)}) : (reg63[(3'h4):(3'h4)] ?
                          reg43 : reg74)) ?
                  ((reg1281[(5'h13):(1'h0)] - (reg44 ? wire1260 : reg101)) ?
                      ($signed(forvar1293) ?
                          wire1291 : (reg1281 ?
                              reg16 : reg1266)) : $unsigned((~^reg1221))) : reg1281[(1'h0):(1'h0)]) ?
              (($unsigned(reg105) >>> $signed(reg1213[(1'h0):(1'h0)])) ?
                  reg1229[(1'h0):(1'h0)] : $signed(((wire2 <<< reg1297) ?
                      $unsigned(reg1298) : (reg1225 + reg95)))) : ((reg1281[(4'hd):(4'hd)] ?
                  (~&(reg70 ?
                      wire1260 : reg1292)) : ({reg1245} << reg16[(2'h2):(2'h2)])) <<< (~(-(&(8'ha3)))))))
            begin
              reg1300 <= $unsigned({$unsigned((reg75[(3'h7):(2'h2)] ?
                      (~^reg1259) : reg1298[(1'h1):(1'h1)]))});
            end
          else
            begin
              reg1301 = (((reg1223 && (^$signed(reg17))) ?
                  (|reg1276[(4'h9):(3'h7)]) : (reg116 ?
                      $unsigned(((8'hbe) ?
                          reg116 : reg1269)) : wire120[(5'h10):(2'h3)])) ~^ $unsigned({reg1213[(1'h0):(1'h0)],
                  ((^reg14) ? $signed(reg1240) : (!reg109))}));
              reg1302 = (7'h44);
              reg1303 <= $signed($unsigned($unsigned(({reg95} ?
                  reg1216 : $signed(reg1213)))));
            end
        end
      else
        begin
          reg1300 <= (&reg99);
          if (forvar1292[(3'h6):(3'h4)])
            begin
              reg1303 <= ((~reg1254) ?
                  ((((reg1263 ? reg85 : reg55) ? (~&reg101) : (~reg40)) ?
                      (&reg45[(4'ha):(4'ha)]) : reg1300[(4'ha):(2'h3)]) == $unsigned((7'h4a))) : reg108[(2'h2):(1'h0)]);
              reg1304 = $unsigned({{$unsigned(reg1277),
                      $unsigned((-reg1267))}});
              reg1305 <= {$unsigned((~&$signed((^reg1298))))};
              reg1306 <= $signed($unsigned($signed(reg1297)));
              reg1307 <= ($unsigned($unsigned(((reg1286 ?
                  wire4 : reg1305) ~^ $signed(reg1263)))) & (|({$unsigned(reg1271),
                      (reg1281 ? reg37 : reg87)} ?
                  (reg37 > $signed((8'ha8))) : ($unsigned(reg1224) & reg108[(1'h0):(1'h0)]))));
            end
          else
            begin
              reg1303 <= ((!wire1290) >>> $unsigned($signed($signed((reg1306 ?
                  reg69 : (8'ha8))))));
              reg1305 <= $unsigned($signed($signed(((reg63 && reg83) ?
                  $unsigned((8'had)) : {reg26, (8'h9e)}))));
              reg1306 <= $unsigned(reg1297[(2'h2):(2'h2)]);
            end
          for (forvar1308 = (1'h0); (forvar1308 < (2'h2)); forvar1308 = (forvar1308 + (1'h1)))
            begin
              reg1309 = reg42;
              reg1310 = $unsigned((~&{reg1271}));
              reg1311 <= reg83[(1'h1):(1'h0)];
              reg1312 = reg82[(4'hb):(4'h9)];
            end
          for (forvar1313 = (1'h0); (forvar1313 < (2'h3)); forvar1313 = (forvar1313 + (1'h1)))
            begin
              reg1314 <= reg1306;
              reg1315 = reg1235;
              reg1316 = reg116;
              reg1317 = ((~&{reg15}) ?
                  ($unsigned((~^reg109)) ?
                      $unsigned((!reg1311)) : ((reg57[(4'h9):(4'h8)] ?
                              (reg1309 ^ reg1310) : (wire1260 <= reg1266)) ?
                          ($unsigned((8'hb6)) * wire1261) : $signed((reg1314 ?
                              reg108 : reg1240)))) : $signed(((-$unsigned(reg1228)) != {$signed((7'h46)),
                      reg1227[(2'h3):(2'h3)]})));
              reg1318 = $unsigned($signed($signed(reg1302)));
            end
          for (forvar1319 = (1'h0); (forvar1319 < (3'h4)); forvar1319 = (forvar1319 + (1'h1)))
            begin
              reg1320 <= $signed((reg63 ? reg95 : reg1301));
              reg1321 <= (~&{((^~(reg31 <= reg1316)) <= reg1223[(4'h9):(3'h4)]),
                  (reg41 ?
                      (~|reg83[(1'h0):(1'h0)]) : $signed((reg17 >= (7'h46))))});
            end
        end
      if (reg72[(4'he):(3'h6)])
        begin
          if (((-reg1307[(4'h8):(2'h3)]) ^~ ((({wire1,
                  wire2} * $unsigned(reg22)) ?
              ($signed(reg70) && $unsigned(reg1315)) : reg99[(4'h8):(4'h8)]) ~^ $signed(($unsigned((8'ha2)) << $unsigned(reg34))))))
            begin
              reg1322 = (($signed(reg1246[(1'h1):(1'h1)]) ^ (((wire4 * (8'ha4)) ?
                      {reg1259} : reg15[(4'hb):(3'h7)]) ?
                  (~(reg14 && reg15)) : reg1302[(4'h9):(1'h0)])) * reg40);
              reg1323 <= (7'h46);
              reg1324 = ({$unsigned($signed((!reg1317))),
                      reg1229[(3'h4):(1'h1)]} ?
                  (reg1309 ?
                      {$unsigned({reg1310})} : $signed({$signed(reg108)})) : $unsigned((&{reg93[(4'hb):(4'hb)]})));
              reg1325 = (~|$unsigned($unsigned($signed((~&reg1277)))));
              reg1326 = (^~wire1260[(4'h9):(3'h5)]);
            end
          else
            begin
              reg1323 <= (reg1225 ?
                  (reg1317 <= (wire1290[(2'h3):(2'h3)] & (reg1317[(1'h0):(1'h0)] ?
                      (+reg1324) : (^reg111)))) : ($signed(($signed(reg97) && (reg1276 ?
                          reg31 : (8'ha4)))) ?
                      (((&reg1318) ?
                          (reg1325 ?
                              reg31 : wire1) : $unsigned(reg1309)) > $signed((~reg87))) : ((&(reg1317 == (8'ha1))) ?
                          reg1242[(4'ha):(3'h7)] : {{(7'h47)}})));
              reg1324 = (~|$unsigned((~reg101)));
              reg1325 = ((reg89 ?
                  ((&(^wire120)) * (&{reg1271,
                      wire1290})) : reg1302) <= (reg1323[(3'h7):(1'h0)] << (&((-reg1322) ?
                  (reg1304 + wire4) : reg1325[(2'h3):(1'h0)]))));
              reg1327 <= $signed($unsigned($signed(reg105[(3'h7):(2'h2)])));
            end
          if ((reg1263[(2'h2):(1'h0)] ?
              ({$signed($signed(wire1261))} >= $unsigned(($signed(reg1235) ?
                  {reg1235,
                      reg1233} : (wire120 != reg1298)))) : $unsigned($unsigned(((wire3 ?
                  reg81 : reg91) != $unsigned(reg16))))))
            begin
              reg1328 = $signed(reg1296);
              reg1329 = $unsigned(reg55[(5'h14):(1'h0)]);
              reg1330 <= ($unsigned($signed((8'hb9))) <= reg1296);
              reg1331 <= (!reg55[(4'h9):(1'h1)]);
              reg1332 <= {reg1327[(2'h2):(1'h1)],
                  $signed($signed(((reg100 ? reg1315 : wire4) ?
                      (reg14 > wire1211) : (reg1223 << reg99))))};
            end
          else
            begin
              reg1330 <= (-$unsigned($unsigned(((~^reg1307) > $signed(reg1254)))));
              reg1331 <= (^~$unsigned(reg70[(1'h1):(1'h0)]));
              reg1332 <= reg49;
              reg1333 = $signed(reg1271);
              reg1334 <= wire1291;
            end
        end
      else
        begin
          reg1322 = (&reg1311);
          if ((reg1298[(3'h4):(2'h3)] ?
              $unsigned((!$signed((reg82 >= reg1281)))) : reg1298))
            begin
              reg1323 <= (+{$signed(wire1), wire1290[(3'h6):(2'h2)]});
              reg1327 <= ((!reg1304) >> {reg1240[(4'h8):(1'h1)]});
              reg1330 <= reg74;
            end
          else
            begin
              reg1323 <= reg1227[(3'h5):(2'h2)];
              reg1324 = reg1320;
              reg1325 = reg1311;
              reg1326 = ({reg1233, reg97[(2'h2):(1'h0)]} ?
                  wire1260 : {($signed((reg1305 ? forvar1293 : (8'ha2))) ?
                          (7'h47) : $unsigned($unsigned(reg1242)))});
              reg1328 = $signed(reg1306[(4'he):(3'h4)]);
            end
        end
    end
  assign wire1335 = (((reg26[(4'h9):(3'h5)] ?
                            ($unsigned((8'hb2)) <<< (+reg1234)) : $unsigned((reg1277 ?
                                reg27 : reg1330))) ?
                        (reg67[(3'h6):(1'h1)] ?
                            $unsigned($unsigned(reg55)) : $unsigned((reg109 + reg93))) : ({(wire4 & wire1),
                                reg101} ?
                            (^reg83) : reg81)) + (&({(reg1224 < (8'hbc))} + (!(~^reg99)))));
  assign wire1336 = (reg1334 ?
                        ((~|(|$unsigned(reg1300))) ?
                            $unsigned($unsigned(((8'hbf) ?
                                reg31 : reg108))) : reg1320[(4'ha):(1'h1)]) : {(|$unsigned({reg1276})),
                            reg72[(5'h12):(5'h10)]});
  always
    @(posedge clk) begin
      reg1337 <= reg108;
    end
  always
    @(posedge clk) begin
      reg1338 = reg1296;
      reg1339 = reg1320;
      reg1340 = (reg21[(4'h9):(4'h9)] ?
          (|(reg1216[(2'h3):(1'h0)] ^~ $signed((~(8'ha4))))) : $unsigned((wire1335 == {$signed(reg1223),
              $unsigned(reg11)})));
      reg1341 <= $unsigned(reg1331[(1'h0):(1'h0)]);
    end
  assign wire1342 = $signed(wire0);
  always
    @(posedge clk) begin
      if (((7'h41) + $unsigned((8'hb8))))
        begin
          for (forvar1343 = (1'h0); (forvar1343 < (1'h1)); forvar1343 = (forvar1343 + (1'h1)))
            begin
              reg1344 <= reg37[(2'h2):(2'h2)];
              reg1345 = $unsigned($signed((&reg1281[(4'hf):(4'hf)])));
              reg1346 = $signed($unsigned($signed(reg1323[(2'h3):(1'h0)])));
              reg1347 <= $signed(reg104);
              reg1348 <= (^~($signed((reg1321[(5'h15):(5'h11)] ?
                      {reg111, (8'hb8)} : reg1337)) ?
                  ({(wire1290 ? reg1306 : reg108), wire3[(1'h1):(1'h1)]} ?
                      reg1276 : reg116[(3'h6):(3'h5)]) : $signed((^~(wire1 ?
                      wire1211 : reg1225)))));
            end
        end
      else
        begin
          reg1343 = $signed((wire1342[(2'h3):(1'h0)] ?
              {(reg104[(3'h6):(1'h1)] || $signed(reg1246))} : ($unsigned({wire1260}) ?
                  (~(8'hb4)) : (~^((8'ha2) ? reg1331 : reg1263)))));
          reg1345 = $unsigned(reg1286[(2'h3):(1'h1)]);
        end
      for (forvar1349 = (1'h0); (forvar1349 < (2'h3)); forvar1349 = (forvar1349 + (1'h1)))
        begin
          reg1350 <= (+$unsigned(reg1343));
        end
    end
  always
    @(posedge clk) begin
      if (reg17)
        begin
          reg1351 <= reg1255[(3'h7):(2'h2)];
          for (forvar1352 = (1'h0); (forvar1352 < (2'h2)); forvar1352 = (forvar1352 + (1'h1)))
            begin
              reg1353 = {reg108, $signed(reg11[(5'h17):(3'h6)])};
              reg1354 <= ($unsigned(((^~reg87[(2'h2):(1'h1)]) ?
                  ((reg1254 ? reg1242 : wire1) ?
                      (reg1274 >>> (8'ha7)) : $unsigned(reg1303)) : reg1234)) * (8'haa));
            end
        end
      else
        begin
          reg1352 = (($signed(reg1242[(4'ha):(2'h2)]) * reg43[(3'h4):(3'h4)]) < (($signed($unsigned(wire1261)) ?
                  reg1303[(3'h6):(2'h2)] : $unsigned((-reg42))) ?
              (!(((8'hbb) ? reg110 : reg55) ?
                  (reg1337 ? (8'h9e) : reg116) : ((8'hb2) ?
                      reg1228 : forvar1352))) : $unsigned($signed((reg89 ?
                  wire1291 : (8'haf))))));
          reg1353 = reg1276;
          for (forvar1354 = (1'h0); (forvar1354 < (3'h4)); forvar1354 = (forvar1354 + (1'h1)))
            begin
              reg1355 <= reg74;
              reg1356 <= ($unsigned(reg93) - reg70);
              reg1357 = (&{$unsigned($unsigned((~&forvar1354))),
                  reg105[(4'hd):(4'hc)]});
              reg1358 = reg87;
              reg1359 = reg34;
            end
        end
      for (forvar1360 = (1'h0); (forvar1360 < (3'h4)); forvar1360 = (forvar1360 + (1'h1)))
        begin
          reg1361 = ((~|$unsigned(((8'hbd) || $signed(wire1342)))) ?
              reg1314[(2'h3):(1'h1)] : reg1327[(4'hd):(4'hc)]);
          for (forvar1362 = (1'h0); (forvar1362 < (2'h3)); forvar1362 = (forvar1362 + (1'h1)))
            begin
              reg1363 = wire1290;
              reg1364 = (-reg1358);
              reg1365 <= {reg81[(3'h5):(1'h0)]};
              reg1366 = reg87[(3'h5):(1'h0)];
              reg1367 = ((reg101[(4'hf):(3'h6)] ?
                      ((reg1352 ?
                          $signed(reg1348) : {reg13,
                              wire1336}) ^~ $unsigned((~&reg83))) : (|reg1271[(1'h0):(1'h0)])) ?
                  reg1311[(2'h2):(1'h1)] : $unsigned($signed((&$unsigned(reg1331)))));
            end
        end
      if ($signed(({reg69[(4'h8):(2'h2)],
          (reg1305[(1'h1):(1'h0)] ?
              $unsigned(reg1347) : reg1269[(3'h5):(1'h1)])} * $unsigned($signed((-wire4))))))
        begin
          if ((~reg81))
            begin
              reg1368 <= $signed({(^~(~^$unsigned(reg108))), reg1223});
              reg1369 = (({reg1356[(2'h2):(1'h0)]} < $signed($signed($unsigned(reg1278)))) ?
                  {reg1229} : reg1359);
              reg1370 <= {$signed(((!$unsigned(reg1267)) ?
                      reg1235 : $signed($signed(reg26))))};
              reg1371 = $signed(reg15);
              reg1372 <= (~^reg1263);
            end
          else
            begin
              reg1368 <= ($unsigned(reg111) > (wire1342 ^ ($signed({reg75}) != (^~reg1221))));
              reg1369 = (~&(^($unsigned({reg1292}) ^~ (reg1334 == $signed(reg1227)))));
              reg1371 = (({{(-reg83), $signed(reg1278)}} ?
                  forvar1354 : reg97) | (~((^~reg1321) ?
                  (7'h47) : ({reg1225} ?
                      $unsigned(reg1296) : (reg37 ? forvar1360 : reg87)))));
              reg1372 <= {{{(reg43 ? $signed(reg1259) : reg16)},
                      ($unsigned($signed(reg110)) ?
                          ($unsigned(wire1261) | (^~reg1369)) : reg99[(2'h3):(2'h3)])}};
            end
          if (((^reg1281[(2'h3):(1'h0)]) ?
              reg1303[(4'h9):(3'h6)] : $signed($unsigned(reg1259[(2'h2):(1'h0)]))))
            begin
              reg1373 = (|reg45[(3'h7):(3'h6)]);
              reg1374 <= ($signed($unsigned($signed((reg1266 << reg43)))) ?
                  $unsigned(((~^$signed((8'hbe))) > (reg81 ?
                      (reg1228 ?
                          (8'haf) : (8'hae)) : $unsigned(wire3)))) : {$signed(((reg1295 * reg1246) - reg1259))});
              reg1375 <= $signed($signed((({reg1277,
                  forvar1362} >= $unsigned(reg1320)) < $signed(reg16[(5'h16):(5'h11)]))));
              reg1376 <= ((~&reg1307[(4'hc):(4'ha)]) ?
                  $signed($signed($signed($unsigned(reg1350)))) : (~&(~|$signed($signed(reg1334)))));
            end
          else
            begin
              reg1374 <= ((reg13[(3'h7):(2'h2)] - ($signed(reg1330[(3'h5):(2'h2)]) ^ $signed((reg89 ?
                      reg82 : (8'ha9))))) ?
                  $unsigned((^~{reg1242[(3'h7):(3'h6)]})) : ($signed($unsigned($unsigned(reg1341))) ?
                      reg1365[(4'hf):(4'h9)] : $unsigned($unsigned(reg31))));
              reg1375 <= $unsigned((reg1296[(3'h5):(2'h2)] | (+((reg1281 | forvar1354) > (reg1361 ?
                  reg1327 : reg1222)))));
            end
          if ($unsigned((8'hb2)))
            begin
              reg1377 = $signed((^~$unsigned($signed(reg1366))));
              reg1378 <= $signed(((((reg1366 ? reg97 : (8'hb6)) ?
                      (reg49 ? reg31 : (8'hb7)) : $signed(reg1233)) ?
                  ((reg21 ? reg1221 : reg31) ?
                      $signed(reg1224) : $unsigned((8'hb8))) : (reg70 > (reg1229 ?
                      reg108 : reg55))) ^~ $signed($unsigned((~^reg26)))));
              reg1379 <= ((~|((~|(8'hbd)) ?
                  reg57 : $unsigned($unsigned((8'h9c))))) <= $unsigned($unsigned(($unsigned(reg72) & $unsigned(reg17)))));
              reg1380 = (~{((-(!(8'hb0))) <<< {$signed(reg82)})});
            end
          else
            begin
              reg1378 <= ((~(reg104[(3'h6):(3'h6)] ?
                      (^~(-(8'ha0))) : (reg1373 ?
                          ((7'h47) != (8'h9f)) : reg1254[(2'h3):(2'h3)]))) ?
                  (($unsigned(reg105[(3'h6):(2'h2)]) ?
                          $unsigned(reg1263) : $unsigned((reg55 ?
                              reg1377 : reg1233))) ?
                      reg1246[(4'hc):(3'h4)] : reg1334) : reg1295[(1'h0):(1'h0)]);
              reg1379 <= (+reg1364);
              reg1380 = ((reg1295[(4'hc):(4'hb)] ?
                  reg1300 : reg1240) & reg1331);
              reg1381 = (((^{reg1355[(4'h8):(2'h3)]}) ^ reg87) ?
                  reg1380[(4'h9):(4'h8)] : ((reg1372[(4'ha):(3'h4)] && $unsigned($signed(reg1341))) ?
                      ($unsigned($unsigned((8'haf))) <<< reg83) : reg1277));
              reg1382 <= $signed(((8'ha3) > $signed((&reg1377[(4'hd):(4'hb)]))));
            end
          reg1383 = $signed(wire2[(4'ha):(2'h3)]);
        end
      else
        begin
          for (forvar1368 = (1'h0); (forvar1368 < (1'h1)); forvar1368 = (forvar1368 + (1'h1)))
            begin
              reg1369 = $signed(reg1352[(4'hc):(1'h1)]);
            end
          reg1370 <= (reg1242[(3'h7):(3'h7)] ?
              (&$unsigned(reg41[(4'hd):(4'hc)])) : $unsigned((!({reg1222} ?
                  ((8'haa) >> reg1276) : (^~reg1350)))));
          reg1372 <= ($unsigned(reg69[(3'h6):(3'h6)]) ?
              (wire2[(4'h9):(3'h6)] ?
                  {(|$signed(reg55))} : $unsigned({((8'ha3) ?
                          (8'hbe) : reg1266)})) : $signed(wire120));
          for (forvar1373 = (1'h0); (forvar1373 < (1'h1)); forvar1373 = (forvar1373 + (1'h1)))
            begin
              reg1374 <= reg55;
              reg1375 <= ((((reg81 > $unsigned((8'hb3))) * {$signed(reg1292)}) ?
                  (&$signed((reg1296 ?
                      (8'ha7) : (7'h46)))) : reg1368[(4'hb):(3'h4)]) || (!reg1327[(3'h5):(2'h2)]));
              reg1376 <= ((($signed((reg109 ?
                      reg1359 : wire1336)) ^ ($unsigned(reg34) ^~ wire0[(4'he):(2'h3)])) ?
                  ((!reg57) ?
                      $unsigned($unsigned(reg1292)) : $signed(reg37)) : ((8'h9e) ?
                      ($unsigned(reg75) ?
                          reg11[(5'h11):(5'h10)] : $signed(reg1376)) : ($signed(reg1307) >= reg87))) + (reg1383 ?
                  $signed(reg1303) : {(reg1303[(4'h8):(3'h5)] & ((8'hba) ?
                          reg91 : (8'hb6)))}));
              reg1378 <= ((reg16[(4'hc):(2'h3)] ?
                  ($signed((reg1366 - (8'hac))) ?
                      $signed((reg1224 >> forvar1354)) : (reg1296 ?
                          (reg55 + reg1369) : reg1372)) : ($unsigned(reg108) * reg1379[(4'ha):(1'h0)])) != (+(^~reg1353)));
              reg1379 <= (8'ha1);
            end
        end
      reg1384 <= (reg1225 & $signed(forvar1362[(4'h8):(3'h5)]));
      for (forvar1385 = (1'h0); (forvar1385 < (1'h1)); forvar1385 = (forvar1385 + (1'h1)))
        begin
          reg1386 = $signed($unsigned((&wire0[(4'ha):(2'h2)])));
          reg1387 <= reg1327;
        end
    end
  assign wire1388 = reg67[(4'h8):(3'h5)];
  assign wire1389 = $signed((^$signed(($signed(reg109) || reg1245[(4'ha):(3'h5)]))));
  always
    @(posedge clk) begin
      reg1390 = reg1269;
      reg1391 = ((+{((~|reg1271) ? (reg1376 ? reg1379 : reg1242) : reg1331)}) ?
          (reg1372 | $unsigned($signed(reg1254[(3'h4):(1'h0)]))) : (reg1374 >> $unsigned((&$unsigned(reg40)))));
      reg1392 <= (((~&($signed((8'haa)) == ((8'hb1) < reg1368))) ?
          wire1336[(1'h1):(1'h0)] : reg1384) ^~ ($unsigned(((^reg1351) && (reg1245 << reg1314))) ?
          ($signed(reg1277[(2'h2):(1'h1)]) > (|reg1295[(4'hb):(3'h5)])) : $unsigned(reg1379)));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module121
#(parameter param1210 = (((+({(8'hb9)} <<< ((8'hb3) ? (8'hb6) : (8'ha9)))) < ((~&((8'ha9) ? (7'h46) : (8'hb1))) + ({(8'hb8), (8'hb8)} != ((8'ha6) < (8'hb0))))) - ((^~(!((8'ha0) >>> (7'h43)))) ? (^~(~&((7'h4a) | (8'hae)))) : ((((8'hb3) - (8'ha9)) ? ((8'hb7) && (7'h41)) : ((8'had) ? (7'h42) : (8'ha2))) ? (|((8'hb6) >> (8'hac))) : (+((8'hb1) ? (8'hb7) : (7'h48)))))))
(y, clk, wire122, wire123, wire124, wire125);
  output wire [(32'h4e7):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(5'h16):(1'h0)] wire122;
  input wire signed [(4'hd):(1'h0)] wire123;
  input wire signed [(3'h5):(1'h0)] wire124;
  input wire signed [(3'h5):(1'h0)] wire125;
  wire signed [(5'h15):(1'h0)] wire126;
  wire [(5'h10):(1'h0)] wire150;
  wire [(3'h5):(1'h0)] wire151;
  wire [(5'h17):(1'h0)] wire194;
  wire [(5'h15):(1'h0)] wire580;
  wire signed [(4'ha):(1'h0)] wire582;
  wire [(3'h5):(1'h0)] wire583;
  wire [(5'h16):(1'h0)] wire1203;
  wire signed [(3'h7):(1'h0)] wire1205;
  wire [(5'h15):(1'h0)] wire1206;
  wire [(4'hb):(1'h0)] wire1207;
  wire [(4'hf):(1'h0)] wire1208;
  reg [(4'h9):(1'h0)] reg596 = (1'h0);
  reg [(5'h15):(1'h0)] reg593 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg589 = (1'h0);
  reg [(5'h11):(1'h0)] reg588 = (1'h0);
  reg [(5'h16):(1'h0)] reg585 = (1'h0);
  reg [(5'h15):(1'h0)] reg193 = (1'h0);
  reg [(5'h16):(1'h0)] reg187 = (1'h0);
  reg [(4'hb):(1'h0)] reg191 = (1'h0);
  reg [(5'h14):(1'h0)] reg190 = (1'h0);
  reg [(5'h11):(1'h0)] reg185 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg182 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg178 = (1'h0);
  reg [(3'h5):(1'h0)] reg177 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg170 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg167 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg163 = (1'h0);
  reg [(5'h10):(1'h0)] reg162 = (1'h0);
  reg [(4'hc):(1'h0)] reg161 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg159 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg158 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg156 = (1'h0);
  reg [(3'h6):(1'h0)] reg155 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg153 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg152 = (1'h0);
  reg [(3'h6):(1'h0)] reg144 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg143 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg142 = (1'h0);
  reg [(5'h17):(1'h0)] reg140 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg138 = (1'h0);
  reg [(4'h8):(1'h0)] reg137 = (1'h0);
  reg [(4'hc):(1'h0)] reg135 = (1'h0);
  reg [(5'h15):(1'h0)] reg134 = (1'h0);
  reg [(5'h14):(1'h0)] reg132 = (1'h0);
  reg [(4'h9):(1'h0)] reg130 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg128 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg127 = (1'h0);
  reg [(5'h10):(1'h0)] reg597 = (1'h0);
  reg [(5'h10):(1'h0)] reg595 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg594 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg592 = (1'h0);
  reg [(5'h13):(1'h0)] reg591 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg590 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg587 = (1'h0);
  reg [(4'hb):(1'h0)] reg586 = (1'h0);
  reg [(4'he):(1'h0)] reg584 = (1'h0);
  reg [(5'h10):(1'h0)] reg192 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg189 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg188 = (1'h0);
  reg [(4'hb):(1'h0)] forvar187 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg186 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg184 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg183 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg181 = (1'h0);
  reg [(4'hb):(1'h0)] reg180 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg179 = (1'h0);
  reg signed [(5'h12):(1'h0)] forvar176 = (1'h0);
  reg [(4'h9):(1'h0)] reg175 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg174 = (1'h0);
  reg [(5'h11):(1'h0)] reg173 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar172 = (1'h0);
  reg [(4'hb):(1'h0)] reg171 = (1'h0);
  reg [(4'ha):(1'h0)] reg169 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar168 = (1'h0);
  reg [(4'hb):(1'h0)] forvar166 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar165 = (1'h0);
  reg [(4'he):(1'h0)] reg164 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg160 = (1'h0);
  reg [(5'h13):(1'h0)] reg157 = (1'h0);
  reg signed [(4'he):(1'h0)] reg154 = (1'h0);
  reg [(3'h5):(1'h0)] reg149 = (1'h0);
  reg [(4'hb):(1'h0)] forvar148 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg147 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg146 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg145 = (1'h0);
  reg [(4'hb):(1'h0)] forvar143 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg136 = (1'h0);
  reg [(3'h5):(1'h0)] forvar131 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg141 = (1'h0);
  reg [(4'h9):(1'h0)] reg139 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar136 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg133 = (1'h0);
  reg [(4'he):(1'h0)] reg131 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg129 = (1'h0);
  assign y = {wire126,
                 wire150,
                 wire151,
                 wire194,
                 wire580,
                 wire582,
                 wire583,
                 wire1203,
                 wire1205,
                 wire1206,
                 wire1207,
                 wire1208,
                 reg596,
                 reg593,
                 reg589,
                 reg588,
                 reg585,
                 reg193,
                 reg187,
                 reg191,
                 reg190,
                 reg185,
                 reg182,
                 reg178,
                 reg177,
                 reg170,
                 reg167,
                 reg163,
                 reg162,
                 reg161,
                 reg159,
                 reg158,
                 reg156,
                 reg155,
                 reg153,
                 reg152,
                 reg144,
                 reg143,
                 reg142,
                 reg140,
                 reg138,
                 reg137,
                 reg135,
                 reg134,
                 reg132,
                 reg130,
                 reg128,
                 reg127,
                 reg597,
                 reg595,
                 reg594,
                 reg592,
                 reg591,
                 reg590,
                 reg587,
                 reg586,
                 reg584,
                 reg192,
                 reg189,
                 reg188,
                 forvar187,
                 reg186,
                 reg184,
                 reg183,
                 reg181,
                 reg180,
                 reg179,
                 forvar176,
                 reg175,
                 reg174,
                 reg173,
                 forvar172,
                 reg171,
                 reg169,
                 forvar168,
                 forvar166,
                 forvar165,
                 reg164,
                 reg160,
                 reg157,
                 reg154,
                 reg149,
                 forvar148,
                 reg147,
                 reg146,
                 reg145,
                 forvar143,
                 reg136,
                 forvar131,
                 reg141,
                 reg139,
                 forvar136,
                 reg133,
                 reg131,
                 reg129,
                 (1'h0)};
  assign wire126 = wire123;
  always
    @(posedge clk) begin
      reg127 <= wire126;
    end
  always
    @(posedge clk) begin
      reg128 <= ((($unsigned($signed((8'h9d))) ?
              wire126[(3'h4):(3'h4)] : $unsigned(wire122[(4'h9):(3'h4)])) ?
          $unsigned(((!wire122) == (reg127 ^ wire125))) : ((wire124 < (wire122 ?
                  wire125 : wire126)) ?
              $unsigned($unsigned((7'h4a))) : wire126[(5'h13):(3'h4)])) ^ $signed($signed((|$unsigned(reg127)))));
      reg129 = {{$signed((^(|wire122))), (~&$unsigned($unsigned(reg127)))}};
      reg130 <= $signed($signed($signed($signed((reg129 ? reg129 : wire123)))));
      if ((+{wire122}))
        begin
          if ((~^($signed($signed($signed(wire123))) <= wire122)))
            begin
              reg131 = reg130[(2'h2):(2'h2)];
              reg132 <= $signed($unsigned((($signed(reg128) <<< wire122[(3'h5):(2'h3)]) * $signed((wire122 ?
                  reg127 : wire123)))));
              reg133 = $unsigned(wire125[(3'h5):(2'h2)]);
              reg134 <= (~{((~^$signed(wire125)) < reg133),
                  ($signed($unsigned(reg129)) ?
                      reg130 : ($signed(wire124) <= $unsigned((7'h46))))});
              reg135 <= ((!(8'h9e)) ?
                  ((~wire125[(3'h5):(2'h3)]) ?
                      {reg129[(1'h1):(1'h0)],
                          ((reg132 ?
                              reg128 : wire125) | {reg127})} : $unsigned((reg130[(4'h8):(4'h8)] >= (reg128 ?
                          reg127 : (7'h45))))) : (~(wire125[(2'h2):(1'h1)] <<< $unsigned((wire125 ?
                      wire126 : wire124)))));
            end
          else
            begin
              reg131 = reg130;
              reg132 <= ($signed($unsigned(((8'ha7) ?
                      (^~(8'ha7)) : $unsigned(reg127)))) ?
                  ((7'h49) <= $signed($unsigned($signed(reg134)))) : (($signed(reg128[(4'hf):(4'hd)]) <= $unsigned($signed(reg128))) ?
                      $unsigned($unsigned($unsigned(wire125))) : $unsigned(reg129[(1'h1):(1'h1)])));
              reg134 <= (~|wire124[(2'h2):(1'h0)]);
            end
          for (forvar136 = (1'h0); (forvar136 < (3'h4)); forvar136 = (forvar136 + (1'h1)))
            begin
              reg137 <= reg131[(3'h4):(1'h0)];
              reg138 <= reg130;
            end
          if ($unsigned((+reg127)))
            begin
              reg139 = $unsigned(($signed({(reg130 ? wire123 : wire124),
                  $signed(wire126)}) + $unsigned((reg138[(2'h2):(2'h2)] >> (forvar136 ?
                  forvar136 : wire124)))));
            end
          else
            begin
              reg140 <= reg127;
              reg141 = $signed(reg130);
              reg142 <= forvar136[(1'h0):(1'h0)];
              reg143 <= $unsigned(reg131);
            end
          reg144 <= reg143;
        end
      else
        begin
          for (forvar131 = (1'h0); (forvar131 < (2'h2)); forvar131 = (forvar131 + (1'h1)))
            begin
              reg133 = {(wire126 ?
                      wire122[(5'h14):(4'he)] : reg129[(1'h0):(1'h0)])};
              reg136 = $unsigned(wire126[(5'h14):(3'h4)]);
              reg139 = (8'h9f);
              reg140 <= (reg141[(2'h3):(2'h2)] ^ $signed(reg130));
              reg141 = ((((reg140[(3'h6):(3'h6)] > {reg128}) << $unsigned(reg143)) <<< (($signed((8'hbe)) ?
                      $unsigned(reg143) : reg127[(4'hf):(4'hb)]) ?
                  (^forvar131) : (^~(8'hb4)))) <<< {(reg142 >>> $signed((wire122 ?
                      (7'h40) : reg137)))});
            end
          reg142 <= (reg129[(3'h6):(3'h6)] >= ((+(reg139 + reg141[(2'h2):(2'h2)])) ?
              ((-$unsigned((8'hbc))) | (reg139 ?
                  $signed((8'hb0)) : reg142)) : $unsigned(reg136[(1'h0):(1'h0)])));
          for (forvar143 = (1'h0); (forvar143 < (1'h0)); forvar143 = (forvar143 + (1'h1)))
            begin
              reg145 = ((+$signed(({forvar136} ?
                  (wire125 && reg129) : $signed(reg134)))) >>> $unsigned(reg132));
              reg146 = ({reg127} >> (reg135 ?
                  (wire123[(3'h7):(3'h6)] ?
                      $signed(wire124[(3'h4):(2'h3)]) : $signed({wire125})) : ((|reg136) ^ ($signed(forvar143) ?
                      (^reg140) : reg145[(4'he):(3'h7)]))));
            end
          reg147 = $signed(($signed(reg130[(3'h7):(3'h6)]) ?
              (((reg138 && (8'ha5)) ?
                  (reg138 - forvar131) : (^~reg141)) >>> (+$unsigned(reg143))) : (~reg138[(1'h0):(1'h0)])));
          for (forvar148 = (1'h0); (forvar148 < (3'h4)); forvar148 = (forvar148 + (1'h1)))
            begin
              reg149 = reg130[(4'h8):(3'h4)];
            end
        end
    end
  assign wire150 = reg132[(4'hb):(3'h5)];
  assign wire151 = $signed((($signed((reg130 * reg144)) >> wire124[(3'h4):(1'h0)]) >= (~|(!$signed(reg130)))));
  always
    @(posedge clk) begin
      reg152 <= ((-{(~$signed(reg135)), $unsigned((reg135 << wire126))}) ?
          (^~reg134[(4'h8):(4'h8)]) : {(~&((reg137 ? (8'ha3) : reg130) ?
                  (8'hbe) : (!reg132))),
              $signed($signed((~^wire122)))});
      if (((reg127[(4'hd):(3'h4)] ?
          (reg134[(1'h1):(1'h1)] <<< ((wire150 ?
              reg135 : wire124) + ((8'haa) & wire151))) : reg152[(3'h6):(3'h4)]) & (-($signed((reg140 ?
              reg127 : reg132)) ?
          ($unsigned(reg128) ?
              $signed(reg127) : wire126[(4'he):(1'h0)]) : ((^reg143) ?
              wire124[(1'h1):(1'h0)] : $signed(reg143))))))
        begin
          reg153 <= {(+$unsigned((((8'hac) < (8'ha7)) ?
                  (reg144 >> wire126) : (|reg134))))};
          reg154 = $signed($unsigned(($signed((+reg134)) ?
              reg137[(1'h1):(1'h1)] : ($signed(wire125) & $unsigned(wire151)))));
          reg155 <= (7'h43);
          reg156 <= reg130[(2'h3):(2'h2)];
          if (($signed($signed(({reg132} ?
              (&(8'h9c)) : (wire150 > wire126)))) ~^ $signed($signed($unsigned((reg143 != (8'hab)))))))
            begin
              reg157 = ($signed((+$unsigned({reg152}))) | (~|($signed(reg130[(1'h1):(1'h1)]) >> ({wire124} ?
                  $unsigned(reg132) : $signed(reg156)))));
              reg158 <= (((wire126[(4'ha):(3'h4)] | {reg157[(5'h10):(5'h10)],
                      ((8'hbd) ^ reg137)}) == (^~reg154[(3'h4):(2'h3)])) ?
                  {$signed(reg140), (!reg143[(3'h6):(1'h0)])} : (7'h42));
              reg159 <= {{$unsigned((!$signed(wire126))), reg134}};
            end
          else
            begin
              reg157 = (&wire125);
            end
        end
      else
        begin
          reg153 <= reg127[(4'h9):(4'h9)];
          if ({(~|(~&($signed(reg128) ?
                  wire122[(1'h1):(1'h1)] : (reg128 ^~ wire124))))})
            begin
              reg155 <= ($unsigned(({{reg157, wire124},
                          wire150[(3'h7):(3'h6)]} ?
                      {{reg137},
                          {wire125,
                              wire125}} : (reg153[(2'h2):(1'h0)] != $unsigned(reg140)))) ?
                  (^~$unsigned(wire122[(3'h7):(3'h7)])) : (&$unsigned((reg130[(1'h0):(1'h0)] > (reg137 ?
                      wire125 : wire126)))));
            end
          else
            begin
              reg155 <= (!wire125);
              reg156 <= $signed(reg132[(5'h13):(5'h11)]);
              reg157 = (($signed((~^reg154)) ?
                      ($signed((reg143 | reg158)) ?
                          (reg142 >= wire123) : $signed(reg127[(5'h11):(4'h8)])) : wire122) ?
                  $signed((reg154 ?
                      $signed($unsigned(reg157)) : $signed((-reg128)))) : reg158);
              reg158 <= (8'ha0);
            end
          reg159 <= $unsigned((wire123[(4'h9):(4'h9)] ?
              reg159[(2'h3):(2'h3)] : $unsigned(reg132)));
          if ($unsigned((8'hbf)))
            begin
              reg160 = (reg142 >>> ((((reg132 ? reg156 : reg130) << (reg157 ?
                          reg153 : reg140)) ?
                      (wire123[(3'h4):(1'h1)] ?
                          wire126 : {reg154,
                              (7'h40)}) : $signed(wire124[(1'h0):(1'h0)])) ?
                  $unsigned((|(wire124 ?
                      wire123 : reg156))) : (((^~wire150) >>> (reg134 ~^ wire123)) && ((^~reg127) ~^ (wire122 << wire123)))));
              reg161 <= {{($unsigned((reg130 != reg142)) ?
                          reg158[(5'h10):(4'hb)] : reg143[(3'h5):(2'h2)]),
                      reg135},
                  reg155[(3'h5):(3'h4)]};
              reg162 <= wire124;
              reg163 <= $signed({($unsigned($signed((8'ha3))) <= ($unsigned((8'hb8)) ?
                      reg154 : (8'hb4))),
                  reg132});
              reg164 = ($signed($signed((^~(7'h43)))) || $unsigned((8'h9c)));
            end
          else
            begin
              reg161 <= (~&($signed((reg137[(3'h7):(3'h6)] && (reg144 > (8'hab)))) ?
                  (7'h41) : reg159[(3'h5):(1'h1)]));
              reg164 = (((~&reg137[(2'h2):(2'h2)]) ~^ (^{reg127,
                      (reg159 ? wire122 : wire124)})) ?
                  $signed(reg144) : $signed({($unsigned(reg144) ^~ (reg137 << wire122))}));
            end
        end
      for (forvar165 = (1'h0); (forvar165 < (1'h1)); forvar165 = (forvar165 + (1'h1)))
        begin
          for (forvar166 = (1'h0); (forvar166 < (2'h3)); forvar166 = (forvar166 + (1'h1)))
            begin
              reg167 <= ($signed(reg153[(3'h7):(3'h5)]) ?
                  reg152[(1'h0):(1'h0)] : $unsigned(forvar165[(3'h7):(1'h1)]));
            end
          for (forvar168 = (1'h0); (forvar168 < (3'h4)); forvar168 = (forvar168 + (1'h1)))
            begin
              reg169 = reg154[(3'h5):(3'h4)];
              reg170 <= {$signed((~^((^reg155) ? reg128 : (-reg169))))};
              reg171 = ((reg138 ~^ $unsigned(((reg154 | wire123) ?
                  (reg143 ?
                      reg127 : reg127) : $unsigned(reg160)))) + reg144[(3'h4):(1'h0)]);
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar172 = (1'h0); (forvar172 < (3'h4)); forvar172 = (forvar172 + (1'h1)))
        begin
          reg173 = reg167;
          reg174 = ($signed($unsigned(wire126[(4'ha):(2'h2)])) ?
              (wire122[(4'hf):(1'h1)] ?
                  ((7'h44) ?
                      ($unsigned(wire150) ~^ $signed(wire123)) : wire123) : ((&{reg140,
                          reg132}) ?
                      $unsigned({(8'ha4)}) : $signed((reg153 >>> wire150)))) : (~$unsigned($unsigned($unsigned(forvar172)))));
          reg175 = $signed((((reg163[(2'h2):(1'h1)] == (reg128 < wire126)) ?
                  (7'h44) : (reg132[(5'h12):(4'hb)] ?
                      (!wire151) : {reg174, reg132})) ?
              ($unsigned((|reg142)) ?
                  ((reg130 ? reg144 : wire123) ?
                      (reg161 ?
                          reg128 : wire151) : reg163[(2'h3):(2'h2)]) : $signed($signed(reg163))) : $signed(reg130[(3'h7):(3'h5)])));
          for (forvar176 = (1'h0); (forvar176 < (3'h4)); forvar176 = (forvar176 + (1'h1)))
            begin
              reg177 <= reg137[(3'h6):(1'h1)];
              reg178 <= (~&$unsigned((8'ha7)));
              reg179 = $unsigned((&((~^(wire124 ?
                  wire126 : forvar172)) >= reg161[(4'hb):(3'h5)])));
              reg180 = $signed({($signed($unsigned(reg159)) ?
                      reg138 : ($signed(reg161) ?
                          $unsigned(wire122) : $signed(wire122)))});
              reg181 = (~^reg180[(3'h5):(2'h2)]);
            end
        end
      if (((~&reg152[(5'h10):(4'hf)]) >= ((^$unsigned((reg155 * reg134))) ?
          ($signed({(8'ha4),
              reg135}) != ((reg135 & reg158) + reg161[(2'h3):(1'h1)])) : (8'hb1))))
        begin
          if ((~^(8'hb6)))
            begin
              reg182 <= reg181;
              reg183 = {(((8'hac) - forvar172) ^ ($unsigned($unsigned(reg178)) ~^ (|(reg143 ?
                      reg179 : (7'h49)))))};
            end
          else
            begin
              reg183 = reg181;
              reg184 = ($signed(((-((8'hb6) & reg161)) ?
                  wire123 : $signed((reg130 ?
                      reg173 : reg127)))) << $unsigned((((|reg183) <<< reg156) == reg173)));
              reg185 <= $signed($unsigned((wire123 <<< ($signed(reg163) ?
                  wire150[(1'h0):(1'h0)] : $unsigned(reg128)))));
              reg186 = ((({{reg179}, (wire151 <= (8'ha5))} ?
                      ((reg142 >>> reg153) ?
                          (reg138 ?
                              reg158 : reg128) : reg174[(5'h11):(3'h4)]) : (-$unsigned(forvar176))) + ((&(reg174 & (7'h41))) ?
                      wire123[(3'h7):(2'h3)] : reg155)) ?
                  $signed({$signed(reg178[(4'h9):(4'h9)])}) : reg134[(4'hb):(4'ha)]);
            end
          for (forvar187 = (1'h0); (forvar187 < (3'h4)); forvar187 = (forvar187 + (1'h1)))
            begin
              reg188 = (~reg156[(3'h7):(1'h0)]);
              reg189 = reg179;
              reg190 <= {reg183};
              reg191 <= reg161[(3'h4):(1'h1)];
            end
        end
      else
        begin
          if (reg127[(3'h7):(3'h7)])
            begin
              reg183 = (reg175[(3'h4):(2'h2)] ?
                  (forvar176 ?
                      reg181 : (+$unsigned({reg178,
                          reg188}))) : (~|reg163[(1'h1):(1'h1)]));
              reg185 <= reg189[(3'h5):(3'h5)];
            end
          else
            begin
              reg183 = reg135[(3'h7):(1'h0)];
              reg185 <= (reg179[(1'h0):(1'h0)] ?
                  reg180[(1'h1):(1'h1)] : (~|reg140));
              reg187 <= reg163[(1'h0):(1'h0)];
            end
          if (($signed($unsigned(reg128[(3'h7):(2'h2)])) > $signed((((wire122 ?
              reg167 : wire125) + (reg188 ?
              reg127 : reg163)) * (reg190[(1'h1):(1'h0)] ?
              (8'ha4) : reg190[(5'h14):(5'h12)])))))
            begin
              reg188 = reg184[(2'h2):(1'h1)];
            end
          else
            begin
              reg188 = reg130[(3'h5):(3'h4)];
              reg190 <= reg144;
              reg192 = reg187[(4'hb):(2'h3)];
              reg193 <= reg170[(2'h2):(2'h2)];
            end
        end
    end
  assign wire194 = {wire150, wire126[(1'h0):(1'h0)]};
  module195 #() modinst581 (wire580, clk, reg127, reg190, reg163, reg135);
  assign wire582 = $unsigned(reg191);
  assign wire583 = {reg170[(2'h2):(2'h2)]};
  always
    @(posedge clk) begin
      reg584 = reg191[(3'h4):(2'h3)];
      if ($signed($signed((reg143[(4'h9):(3'h4)] ?
          {((8'ha5) ? reg190 : reg170)} : $signed((~^reg134))))))
        begin
          if ((($signed($unsigned(((8'hb0) != wire194))) ?
              $unsigned(((reg177 ?
                  reg167 : reg167) == (wire123 ^ wire194))) : (8'hb1)) ^~ reg178))
            begin
              reg585 <= $signed(reg144);
            end
          else
            begin
              reg586 = ($signed($unsigned(((8'ha2) * $signed((7'h45))))) ?
                  wire194 : ($signed($unsigned((reg152 | reg187))) & $unsigned($signed((8'hbe)))));
              reg587 = (8'ha8);
              reg588 <= {{{$signed((reg182 < reg185)),
                          {(reg153 + reg162), (~&reg193)}}}};
            end
          reg589 <= $signed($unsigned(reg167[(4'he):(4'he)]));
          if (wire580[(5'h13):(4'h9)])
            begin
              reg590 = $signed((8'h9d));
              reg591 = $signed(wire151);
              reg592 = reg191[(2'h2):(1'h0)];
            end
          else
            begin
              reg590 = $unsigned((reg187[(4'h9):(4'h9)] >= reg584[(1'h1):(1'h1)]));
              reg591 = $unsigned($signed((reg167[(4'h9):(3'h5)] ?
                  reg158 : reg193[(4'hc):(2'h2)])));
              reg592 = $unsigned(reg587[(1'h0):(1'h0)]);
              reg593 <= reg137;
            end
        end
      else
        begin
          reg586 = $unsigned(reg142[(3'h6):(1'h1)]);
          reg587 = reg143;
          reg590 = {$signed(({reg593, $unsigned(reg591)} >>> {(!(7'h46))}))};
          if ($signed($signed((-reg187))))
            begin
              reg591 = ($unsigned(((wire122 ?
                  $unsigned(reg177) : {reg167,
                      reg128}) >= reg178)) == $unsigned($unsigned((|$signed(wire580)))));
              reg593 <= $unsigned($unsigned(reg155[(2'h3):(2'h3)]));
              reg594 = $unsigned((~^reg155));
              reg595 = $signed((+(~reg132)));
            end
          else
            begin
              reg593 <= $unsigned(($unsigned(reg593) ?
                  (~&{$unsigned(reg587)}) : ((~$signed((8'hb9))) | reg135)));
              reg594 = (7'h4a);
              reg595 = (reg159[(3'h6):(3'h5)] ?
                  (8'hb6) : ((+reg162) ?
                      reg190[(4'hd):(4'hd)] : $unsigned(reg590)));
              reg596 <= $signed(wire580);
              reg597 = reg143[(1'h1):(1'h1)];
            end
        end
    end
  module598 #() modinst1204 (wire1203, clk, reg135, reg134, reg158, reg193);
  assign wire1205 = reg593[(4'h9):(1'h1)];
  assign wire1206 = $signed($signed($signed(({reg170} + $signed(wire126)))));
  assign wire1207 = $signed(((((+reg589) ? $unsigned(reg156) : wire1205) ?
                            ($unsigned(reg159) ?
                                reg163 : $unsigned((8'hb7))) : $signed($signed(reg589))) ?
                        (~((wire1205 > wire582) ?
                            (8'hb9) : wire125)) : (^(reg596[(1'h0):(1'h0)] << $unsigned(reg134)))));
  module420 #() modinst1209 (.y(wire1208), .wire425(reg585), .wire422(wire580), .wire421(wire122), .wire424(wire125), .wire423(reg153), .clk(clk));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module598  (y, clk, wire602, wire601, wire600, wire599);
  output wire [(32'h429):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(3'h5):(1'h0)] wire602;
  input wire signed [(3'h6):(1'h0)] wire601;
  input wire [(5'h12):(1'h0)] wire600;
  input wire [(5'h15):(1'h0)] wire599;
  wire [(2'h3):(1'h0)] wire1202;
  wire [(4'hb):(1'h0)] wire960;
  wire signed [(5'h15):(1'h0)] wire641;
  wire signed [(4'hf):(1'h0)] wire640;
  wire [(5'h10):(1'h0)] wire607;
  wire signed [(4'hd):(1'h0)] wire606;
  wire [(4'ha):(1'h0)] wire605;
  wire [(5'h17):(1'h0)] wire604;
  wire signed [(4'hd):(1'h0)] wire1164;
  reg signed [(5'h14):(1'h0)] reg1201 = (1'h0);
  reg [(5'h11):(1'h0)] reg1199 = (1'h0);
  reg [(5'h15):(1'h0)] reg1196 = (1'h0);
  reg [(4'he):(1'h0)] reg1192 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1191 = (1'h0);
  reg [(4'he):(1'h0)] reg1188 = (1'h0);
  reg [(4'hf):(1'h0)] reg1185 = (1'h0);
  reg [(5'h16):(1'h0)] reg1184 = (1'h0);
  reg [(5'h10):(1'h0)] reg1183 = (1'h0);
  reg [(3'h4):(1'h0)] reg1182 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1180 = (1'h0);
  reg [(2'h3):(1'h0)] reg1178 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1176 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1175 = (1'h0);
  reg [(5'h11):(1'h0)] reg1173 = (1'h0);
  reg [(2'h2):(1'h0)] reg1171 = (1'h0);
  reg [(5'h16):(1'h0)] reg1170 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg609 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg611 = (1'h0);
  reg [(3'h5):(1'h0)] reg613 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg617 = (1'h0);
  reg [(4'hd):(1'h0)] reg619 = (1'h0);
  reg [(5'h17):(1'h0)] reg620 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg621 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg624 = (1'h0);
  reg [(5'h17):(1'h0)] reg625 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg627 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg628 = (1'h0);
  reg [(2'h3):(1'h0)] reg629 = (1'h0);
  reg [(4'ha):(1'h0)] reg633 = (1'h0);
  reg [(5'h17):(1'h0)] reg634 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg636 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1200 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1198 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar1197 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1195 = (1'h0);
  reg [(5'h13):(1'h0)] reg1194 = (1'h0);
  reg [(5'h17):(1'h0)] forvar1193 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1190 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1186 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1189 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1187 = (1'h0);
  reg [(4'ha):(1'h0)] forvar1186 = (1'h0);
  reg [(3'h6):(1'h0)] reg1181 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1179 = (1'h0);
  reg [(5'h14):(1'h0)] forvar1175 = (1'h0);
  reg [(4'h9):(1'h0)] reg1177 = (1'h0);
  reg [(5'h16):(1'h0)] reg1174 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1172 = (1'h0);
  reg [(5'h17):(1'h0)] reg1169 = (1'h0);
  reg [(2'h2):(1'h0)] reg1168 = (1'h0);
  reg [(3'h7):(1'h0)] reg1167 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar1166 = (1'h0);
  reg [(2'h2):(1'h0)] reg642 = (1'h0);
  reg [(5'h10):(1'h0)] reg639 = (1'h0);
  reg [(5'h16):(1'h0)] reg638 = (1'h0);
  reg [(5'h10):(1'h0)] reg637 = (1'h0);
  reg [(4'h8):(1'h0)] reg635 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg632 = (1'h0);
  reg [(5'h15):(1'h0)] reg631 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg630 = (1'h0);
  reg [(3'h7):(1'h0)] reg626 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg623 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar622 = (1'h0);
  reg [(5'h13):(1'h0)] reg618 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg616 = (1'h0);
  reg [(4'hd):(1'h0)] reg615 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg614 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg612 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar610 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg608 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg603 = (1'h0);
  assign y = {wire1202,
                 wire960,
                 wire641,
                 wire640,
                 wire607,
                 wire606,
                 wire605,
                 wire604,
                 wire1164,
                 reg1201,
                 reg1199,
                 reg1196,
                 reg1192,
                 reg1191,
                 reg1188,
                 reg1185,
                 reg1184,
                 reg1183,
                 reg1182,
                 reg1180,
                 reg1178,
                 reg1176,
                 reg1175,
                 reg1173,
                 reg1171,
                 reg1170,
                 reg609,
                 reg611,
                 reg613,
                 reg617,
                 reg619,
                 reg620,
                 reg621,
                 reg624,
                 reg625,
                 reg627,
                 reg628,
                 reg629,
                 reg633,
                 reg634,
                 reg636,
                 reg1200,
                 reg1198,
                 forvar1197,
                 reg1195,
                 reg1194,
                 forvar1193,
                 reg1190,
                 reg1186,
                 reg1189,
                 reg1187,
                 forvar1186,
                 reg1181,
                 reg1179,
                 forvar1175,
                 reg1177,
                 reg1174,
                 reg1172,
                 reg1169,
                 reg1168,
                 reg1167,
                 forvar1166,
                 reg642,
                 reg639,
                 reg638,
                 reg637,
                 reg635,
                 reg632,
                 reg631,
                 reg630,
                 reg626,
                 reg623,
                 forvar622,
                 reg618,
                 reg616,
                 reg615,
                 reg614,
                 reg612,
                 forvar610,
                 reg608,
                 reg603,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg603 = wire601;
    end
  assign wire604 = {(+(~wire600)),
                       (wire601[(2'h3):(1'h0)] || ($signed($unsigned(wire599)) * $signed(wire601)))};
  assign wire605 = $unsigned((~{((^~wire602) >> $unsigned(wire600)),
                       ((wire602 ? wire602 : wire599) ?
                           ((8'ha6) ?
                               wire601 : wire600) : wire602[(2'h2):(2'h2)])}));
  assign wire606 = $signed({(((7'h47) ?
                           $unsigned(wire601) : (~|wire605)) == wire602[(3'h5):(1'h0)]),
                       wire599});
  assign wire607 = $signed(wire606);
  always
    @(posedge clk) begin
      reg608 = ($signed(wire600[(4'ha):(4'ha)]) <= (~|(((wire607 ?
              wire601 : wire602) <<< $unsigned(wire605)) ?
          (wire604 | (-wire605)) : $signed((wire605 >= wire601)))));
      reg609 <= wire601[(3'h5):(2'h3)];
      for (forvar610 = (1'h0); (forvar610 < (3'h4)); forvar610 = (forvar610 + (1'h1)))
        begin
          if ((((&($unsigned(wire599) | (&wire605))) ?
              ((~((8'ha1) ? forvar610 : forvar610)) >> ({wire607} ?
                  $signed(wire605) : (8'h9c))) : wire601) ^ (($unsigned((8'hb4)) || $unsigned((^wire604))) ?
              wire602[(2'h2):(2'h2)] : (({wire604,
                  wire599} - wire599) != (+wire606)))))
            begin
              reg611 <= {({((wire605 ^ wire604) || (reg609 ?
                          wire602 : (7'h49))),
                      {(wire604 ? wire599 : (8'hab)),
                          $signed(reg609)}} ^~ {((wire607 & (7'h48)) * $signed(wire605)),
                      (8'h9d)})};
              reg612 = (~((&(wire602[(1'h1):(1'h1)] | (wire607 ?
                      (8'hb8) : wire604))) ?
                  (^(~^(reg609 + wire607))) : wire602));
              reg613 <= (+$signed(($unsigned(wire607) * ({wire604} ?
                  (8'hb8) : (~wire606)))));
              reg614 = (|reg611[(5'h13):(2'h2)]);
              reg615 = $signed(($signed($signed(wire602[(2'h2):(2'h2)])) ?
                  (($signed(wire606) < (wire602 ?
                      reg608 : wire601)) >> reg608) : ((!(~|wire599)) ?
                      ($signed((8'hb6)) < wire599) : (reg611 ^~ $signed(wire601)))));
            end
          else
            begin
              reg611 <= ($signed(($signed($unsigned((8'ha7))) ?
                  wire602 : $signed(((8'hbe) ~^ wire604)))) >= reg614[(4'h9):(3'h4)]);
              reg612 = $signed(((((reg613 ? reg615 : wire604) ?
                  {reg612,
                      (7'h46)} : (reg608 >> reg614)) * reg613) + (!(wire600[(4'hd):(4'h8)] ?
                  $unsigned((8'hab)) : wire606))));
            end
          reg616 = reg609;
          if ($unsigned(wire604))
            begin
              reg617 <= wire605[(3'h5):(2'h2)];
              reg618 = (+(reg614 ?
                  ((~|$signed(wire605)) >>> ($unsigned(wire605) ?
                      $unsigned(reg615) : wire606[(1'h1):(1'h1)])) : ({$unsigned(wire599)} & wire604)));
            end
          else
            begin
              reg618 = ($signed((~^(!reg613[(2'h3):(1'h0)]))) ?
                  {$signed(reg614[(4'ha):(4'ha)]),
                      $unsigned((((8'hb6) | (8'hb8)) <<< $signed((8'h9d))))} : (wire606 ?
                      reg614[(3'h4):(2'h2)] : reg611));
              reg619 <= (~wire599);
              reg620 <= (&(forvar610 ?
                  reg619[(2'h3):(1'h1)] : $signed($signed(reg619))));
              reg621 <= $signed(reg619[(4'hc):(3'h6)]);
            end
          for (forvar622 = (1'h0); (forvar622 < (2'h2)); forvar622 = (forvar622 + (1'h1)))
            begin
              reg623 = reg615;
            end
        end
      reg624 <= $unsigned((-reg621));
      reg625 <= reg608[(3'h4):(2'h2)];
    end
  always
    @(posedge clk) begin
      if (reg625)
        begin
          if ($unsigned($unsigned(({{reg621}} ^ (!$signed((7'h4a)))))))
            begin
              reg626 = reg617[(4'hb):(3'h4)];
              reg627 <= (+{wire601[(1'h1):(1'h1)],
                  (!((wire599 ? reg621 : wire601) ^ $unsigned(reg609)))});
              reg628 <= wire606[(1'h1):(1'h0)];
              reg629 <= {((|(8'hb0)) ^~ {$unsigned(reg613[(3'h4):(3'h4)])}),
                  $unsigned($unsigned(reg628))};
              reg630 = ($signed(($unsigned(((7'h41) == wire601)) ?
                  reg627 : (wire606 > $signed(wire600)))) >= reg609[(4'hd):(4'hd)]);
            end
          else
            begin
              reg626 = $signed(((~&(~|$signed((7'h41)))) & $signed($signed((reg620 & reg626)))));
              reg630 = reg626;
              reg631 = ($signed((wire601[(1'h1):(1'h1)] | $signed((8'hb8)))) | $unsigned((reg609 ?
                  (&reg611[(5'h10):(3'h5)]) : ({(8'hac)} ?
                      reg629 : $unsigned((8'ha1))))));
              reg632 = reg628;
            end
          reg633 <= reg620;
          reg634 <= reg621;
          if (reg626)
            begin
              reg635 = ($unsigned($unsigned(($unsigned(reg632) && reg632[(4'hd):(4'h8)]))) - $signed(reg627));
              reg636 <= $unsigned({reg625,
                  (reg634[(5'h16):(3'h4)] >= (+(reg609 ? reg617 : reg609)))});
              reg637 = wire599[(3'h5):(2'h2)];
              reg638 = $signed((~((((8'hb9) < (8'hbe)) << $signed(wire606)) ?
                  (|reg626[(3'h5):(1'h1)]) : ((reg633 > wire600) ?
                      (wire607 ? wire605 : wire600) : $unsigned(wire601)))));
            end
          else
            begin
              reg636 <= ((-wire605[(1'h1):(1'h0)]) >>> wire600[(4'he):(4'hc)]);
            end
        end
      else
        begin
          if (reg620)
            begin
              reg627 <= (^~$unsigned((~&reg638)));
              reg630 = wire601[(1'h0):(1'h0)];
              reg633 <= $unsigned($signed(($signed({reg625,
                  reg637}) ~^ $signed(wire601))));
              reg634 <= reg629;
              reg636 <= $signed(reg620[(4'hb):(3'h4)]);
            end
          else
            begin
              reg626 = $unsigned((-$unsigned((!(reg627 | reg628)))));
              reg630 = wire605[(3'h5):(1'h1)];
              reg633 <= $unsigned((reg619 >= (($signed(reg609) <<< reg611) <<< ($unsigned(wire602) >> {(8'hbb)}))));
              reg635 = ($unsigned(wire604[(4'hc):(1'h0)]) ?
                  reg634 : reg621[(3'h7):(3'h7)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg639 = (($unsigned((wire605 ?
              wire607 : (reg625 ? reg619 : wire605))) - reg613[(2'h3):(1'h0)]) ?
          (~reg619[(4'ha):(4'h8)]) : $unsigned((wire600 ?
              (~^(wire607 ? (8'ha5) : reg636)) : reg625[(4'he):(4'hc)])));
    end
  assign wire640 = $signed((7'h44));
  assign wire641 = $unsigned($unsigned(({(~|reg619), reg609[(3'h6):(1'h0)]} ?
                       reg619[(1'h0):(1'h0)] : (|$signed(reg627)))));
  always
    @(posedge clk) begin
      reg642 = wire604[(4'hd):(4'h9)];
    end
  module643 #() modinst961 (wire960, clk, reg627, reg620, reg624, wire641, reg625);
  module962 #() modinst1165 (wire1164, clk, reg628, reg634, reg627, wire604);
  always
    @(posedge clk) begin
      for (forvar1166 = (1'h0); (forvar1166 < (2'h2)); forvar1166 = (forvar1166 + (1'h1)))
        begin
          reg1167 = reg628;
          if ($signed({(wire960 << forvar1166),
              $signed((|(reg613 + wire640)))}))
            begin
              reg1168 = {$signed($signed(reg620)),
                  (((~&$signed(reg633)) >= reg619[(3'h5):(3'h5)]) >> $signed((wire607 ?
                      (wire641 ? wire600 : wire641) : {reg619, reg624})))};
              reg1169 = $signed((-reg1168[(2'h2):(2'h2)]));
            end
          else
            begin
              reg1168 = (($unsigned($unsigned((~forvar1166))) > $signed($unsigned($unsigned(reg613)))) ?
                  wire606[(3'h4):(1'h1)] : ({wire601[(1'h0):(1'h0)]} ?
                      {(reg609[(3'h5):(1'h1)] ? (reg634 + reg633) : {wire641}),
                          reg620[(1'h1):(1'h0)]} : $signed((reg1168 ?
                          (~^wire599) : forvar1166[(4'h9):(4'h8)]))));
              reg1170 <= {(($unsigned($signed(reg1169)) ?
                      wire607 : $signed($unsigned(reg611))) * ($unsigned({reg629,
                          reg619}) ?
                      reg636 : $signed({(8'hba)})))};
              reg1171 <= {reg633[(1'h1):(1'h0)],
                  ((~^reg625[(4'hf):(2'h3)]) ?
                      (+((reg609 >> (7'h49)) ?
                          ((8'ha0) <<< (8'ha9)) : ((8'haa) | wire604))) : $signed((8'hac)))};
              reg1172 = reg625[(4'ha):(2'h2)];
            end
          reg1173 <= (-$signed({(~&wire600[(3'h4):(2'h3)])}));
          reg1174 = (($unsigned(reg619) - reg636[(1'h1):(1'h1)]) ?
              $unsigned(wire640) : ({wire1164[(2'h3):(1'h0)],
                  reg1167} >> wire960[(3'h4):(2'h2)]));
        end
      if ($signed(($unsigned((8'hb4)) - $unsigned(((|(8'haf)) << (+reg633))))))
        begin
          if ((&$signed((reg628 || wire605))))
            begin
              reg1175 <= {(wire605 << reg1174), $unsigned((8'hbe))};
              reg1176 <= (|$signed((8'ha8)));
            end
          else
            begin
              reg1177 = $unsigned($signed((reg636[(3'h5):(2'h3)] ?
                  reg1168[(1'h1):(1'h1)] : $unsigned(forvar1166[(4'hc):(2'h2)]))));
              reg1178 <= ($signed((wire602[(2'h3):(1'h1)] ^~ ((reg1174 ?
                      reg620 : reg620) ?
                  {reg609,
                      (8'ha6)} : reg1172[(4'h9):(3'h5)]))) >> ({{(reg1169 * wire640),
                          (~|reg611)},
                      ((reg1170 <= reg1176) ^ wire641)} ?
                  (^reg1176) : ((reg634[(5'h10):(4'ha)] >= reg1176[(2'h2):(1'h1)]) ?
                      (wire605 <<< (reg1176 == wire605)) : reg636)));
            end
        end
      else
        begin
          for (forvar1175 = (1'h0); (forvar1175 < (3'h4)); forvar1175 = (forvar1175 + (1'h1)))
            begin
              reg1176 <= reg627[(4'h9):(3'h5)];
              reg1177 = (^~(~&$unsigned(reg613[(1'h0):(1'h0)])));
              reg1179 = reg1171[(2'h2):(2'h2)];
              reg1180 <= {reg1178[(1'h0):(1'h0)], (reg1171 < reg619)};
            end
          reg1181 = wire640[(4'h9):(1'h1)];
          reg1182 <= reg1169[(3'h7):(3'h5)];
          reg1183 <= (+wire602[(3'h4):(2'h3)]);
        end
      if (wire640[(2'h3):(1'h0)])
        begin
          reg1184 <= wire1164[(3'h6):(1'h1)];
          reg1185 <= (~|($signed($signed(((8'h9d) ? reg1175 : reg1171))) ?
              ($unsigned($signed(reg609)) != $unsigned((reg633 ?
                  reg627 : (8'hbe)))) : forvar1166[(4'hc):(4'h8)]));
          for (forvar1186 = (1'h0); (forvar1186 < (3'h4)); forvar1186 = (forvar1186 + (1'h1)))
            begin
              reg1187 = {$signed(forvar1175[(3'h6):(2'h3)])};
              reg1188 <= $signed(reg1181);
            end
          reg1189 = (!{reg1174,
              (~|{(reg617 | reg628), wire600[(4'hb):(4'hb)]})});
        end
      else
        begin
          reg1184 <= reg628;
          reg1186 = $unsigned($unsigned(reg617));
          if ((($signed(reg1174[(2'h3):(1'h0)]) ?
                  $unsigned(reg1185) : forvar1166) ?
              (~^$unsigned($unsigned((&reg1183)))) : $signed(reg1174)))
            begin
              reg1187 = (^$signed(reg1173[(3'h4):(1'h0)]));
              reg1188 <= (($unsigned((~^(wire640 | (8'ha8)))) ?
                      $unsigned(($signed(reg625) ?
                          reg1178[(2'h3):(2'h2)] : (wire640 && reg1180))) : ((~&wire601) ?
                          (~^(+reg1176)) : wire960[(1'h1):(1'h1)])) ?
                  reg1180[(3'h5):(1'h1)] : (|$signed((reg1175[(1'h0):(1'h0)] ?
                      (8'hb1) : (8'hbb)))));
              reg1189 = ($unsigned((~|$unsigned((reg1167 >>> (8'hab))))) ?
                  (^~reg625[(5'h12):(4'he)]) : $signed(reg1178));
              reg1190 = (8'had);
            end
          else
            begin
              reg1188 <= (|($unsigned($signed((reg613 ? reg1184 : reg633))) ?
                  (8'hbd) : {($unsigned(wire960) | reg1175),
                      (reg617 <<< $unsigned(reg627))}));
              reg1191 <= reg1185[(1'h0):(1'h0)];
              reg1192 <= ($signed(reg1184) - wire600[(3'h4):(3'h4)]);
            end
        end
      for (forvar1193 = (1'h0); (forvar1193 < (3'h4)); forvar1193 = (forvar1193 + (1'h1)))
        begin
          reg1194 = (forvar1186[(4'h9):(3'h6)] < ((|({(8'haa),
              reg1178} != (8'hbf))) < reg1173));
          reg1195 = (~&$signed(($signed(reg1188) ?
              {$unsigned(reg1189), $unsigned((8'ha9))} : {reg1176})));
          reg1196 <= ((^~reg611[(5'h11):(4'he)]) ~^ ({reg611,
                  (|$unsigned(wire641))} ?
              {wire600[(3'h7):(2'h2)]} : (reg611 ?
                  reg1176 : forvar1193[(5'h16):(1'h1)])));
          for (forvar1197 = (1'h0); (forvar1197 < (2'h2)); forvar1197 = (forvar1197 + (1'h1)))
            begin
              reg1198 = $unsigned(reg1178);
              reg1199 <= (8'h9f);
              reg1200 = (($signed((^~wire601)) ?
                  $signed($unsigned((reg1168 ?
                      reg1172 : reg1174))) : ($signed(reg1171) - reg1167[(3'h6):(3'h6)])) | (wire599[(2'h2):(2'h2)] ?
                  (~&reg627[(3'h4):(2'h2)]) : (+($signed(wire641) ?
                      (~|reg1175) : $signed(wire600)))));
              reg1201 <= ($unsigned((((reg611 ? reg1175 : reg1194) - reg1199) ?
                  $unsigned((8'ha5)) : reg634[(4'h8):(1'h1)])) & wire960);
            end
        end
    end
  assign wire1202 = reg613[(3'h5):(2'h3)];
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module195
#(parameter param579 = (~|(~&((((8'hb9) >>> (8'ha9)) ^ ((8'hb9) >>> (7'h41))) ? (!(|(8'haf))) : (+((8'hb0) && (8'h9f)))))))
(y, clk, wire199, wire198, wire197, wire196);
  output wire [(32'hc1b):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire199;
  input wire [(4'h8):(1'h0)] wire198;
  input wire signed [(5'h18):(1'h0)] wire197;
  input wire [(4'hb):(1'h0)] wire196;
  wire signed [(5'h15):(1'h0)] wire578;
  wire [(3'h7):(1'h0)] wire577;
  wire signed [(3'h6):(1'h0)] wire575;
  wire signed [(2'h3):(1'h0)] wire407;
  wire signed [(4'hd):(1'h0)] wire403;
  wire [(3'h4):(1'h0)] wire402;
  wire signed [(4'ha):(1'h0)] wire379;
  wire [(4'ha):(1'h0)] wire345;
  wire [(5'h11):(1'h0)] wire323;
  wire signed [(2'h2):(1'h0)] wire221;
  wire [(4'hd):(1'h0)] wire200;
  reg signed [(2'h2):(1'h0)] reg203 = (1'h0);
  reg [(4'h9):(1'h0)] reg204 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg205 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg209 = (1'h0);
  reg [(4'hc):(1'h0)] reg210 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg211 = (1'h0);
  reg [(3'h6):(1'h0)] reg213 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg214 = (1'h0);
  reg [(5'h17):(1'h0)] reg217 = (1'h0);
  reg [(4'hc):(1'h0)] reg220 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg225 = (1'h0);
  reg [(5'h16):(1'h0)] reg227 = (1'h0);
  reg [(5'h18):(1'h0)] reg228 = (1'h0);
  reg [(4'hb):(1'h0)] reg230 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg231 = (1'h0);
  reg [(4'hd):(1'h0)] reg232 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg233 = (1'h0);
  reg [(5'h17):(1'h0)] reg235 = (1'h0);
  reg [(5'h13):(1'h0)] reg242 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg244 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg245 = (1'h0);
  reg [(5'h10):(1'h0)] reg247 = (1'h0);
  reg [(5'h16):(1'h0)] reg248 = (1'h0);
  reg [(4'he):(1'h0)] reg249 = (1'h0);
  reg [(4'he):(1'h0)] reg251 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg256 = (1'h0);
  reg [(5'h14):(1'h0)] reg257 = (1'h0);
  reg [(3'h4):(1'h0)] reg258 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg259 = (1'h0);
  reg [(5'h13):(1'h0)] reg260 = (1'h0);
  reg [(2'h2):(1'h0)] reg263 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg264 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg268 = (1'h0);
  reg [(5'h16):(1'h0)] reg271 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg273 = (1'h0);
  reg [(4'h9):(1'h0)] reg276 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg280 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg281 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg283 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg284 = (1'h0);
  reg [(2'h3):(1'h0)] reg286 = (1'h0);
  reg [(5'h18):(1'h0)] reg288 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg291 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg292 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg293 = (1'h0);
  reg [(4'h8):(1'h0)] reg294 = (1'h0);
  reg [(3'h6):(1'h0)] reg299 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg301 = (1'h0);
  reg [(3'h4):(1'h0)] reg308 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg311 = (1'h0);
  reg [(4'hc):(1'h0)] reg313 = (1'h0);
  reg [(4'ha):(1'h0)] reg316 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg318 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg322 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg325 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg326 = (1'h0);
  reg [(5'h16):(1'h0)] reg327 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg328 = (1'h0);
  reg [(2'h2):(1'h0)] reg329 = (1'h0);
  reg [(4'h8):(1'h0)] reg332 = (1'h0);
  reg [(4'ha):(1'h0)] reg333 = (1'h0);
  reg [(5'h14):(1'h0)] reg331 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg334 = (1'h0);
  reg [(5'h16):(1'h0)] reg337 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg339 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg341 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg336 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg342 = (1'h0);
  reg [(4'hf):(1'h0)] reg347 = (1'h0);
  reg [(4'hb):(1'h0)] reg348 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg349 = (1'h0);
  reg [(5'h18):(1'h0)] reg350 = (1'h0);
  reg [(4'hc):(1'h0)] reg351 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg356 = (1'h0);
  reg [(4'he):(1'h0)] reg357 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg359 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg360 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg362 = (1'h0);
  reg [(4'hb):(1'h0)] reg363 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg364 = (1'h0);
  reg [(4'h8):(1'h0)] reg367 = (1'h0);
  reg [(5'h11):(1'h0)] reg369 = (1'h0);
  reg [(5'h14):(1'h0)] reg371 = (1'h0);
  reg [(5'h10):(1'h0)] reg372 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg373 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg377 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg378 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg382 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg385 = (1'h0);
  reg [(5'h11):(1'h0)] reg387 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg384 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg386 = (1'h0);
  reg [(4'hf):(1'h0)] reg391 = (1'h0);
  reg [(5'h12):(1'h0)] reg395 = (1'h0);
  reg [(3'h5):(1'h0)] reg399 = (1'h0);
  reg [(4'hd):(1'h0)] reg400 = (1'h0);
  reg [(5'h17):(1'h0)] reg404 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg406 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg408 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg409 = (1'h0);
  reg [(5'h14):(1'h0)] reg412 = (1'h0);
  reg [(4'he):(1'h0)] reg414 = (1'h0);
  reg [(5'h10):(1'h0)] reg419 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg418 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg417 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg416 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg415 = (1'h0);
  reg [(2'h3):(1'h0)] reg413 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar411 = (1'h0);
  reg [(4'hb):(1'h0)] forvar410 = (1'h0);
  reg [(4'hc):(1'h0)] forvar405 = (1'h0);
  reg [(4'h9):(1'h0)] reg401 = (1'h0);
  reg [(5'h14):(1'h0)] reg398 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar397 = (1'h0);
  reg [(2'h2):(1'h0)] reg396 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg394 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg393 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar392 = (1'h0);
  reg [(5'h17):(1'h0)] forvar390 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg389 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg388 = (1'h0);
  reg [(3'h7):(1'h0)] forvar386 = (1'h0);
  reg [(4'hb):(1'h0)] forvar384 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg383 = (1'h0);
  reg [(5'h14):(1'h0)] reg381 = (1'h0);
  reg [(5'h10):(1'h0)] reg380 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar376 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg375 = (1'h0);
  reg [(5'h16):(1'h0)] reg374 = (1'h0);
  reg [(4'h8):(1'h0)] reg370 = (1'h0);
  reg [(4'hf):(1'h0)] reg368 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg366 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg365 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg361 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg358 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg355 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg354 = (1'h0);
  reg [(4'hd):(1'h0)] reg353 = (1'h0);
  reg [(3'h7):(1'h0)] reg352 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar346 = (1'h0);
  reg [(4'hf):(1'h0)] reg344 = (1'h0);
  reg [(4'hb):(1'h0)] reg343 = (1'h0);
  reg [(5'h13):(1'h0)] reg340 = (1'h0);
  reg [(4'hf):(1'h0)] reg338 = (1'h0);
  reg [(5'h16):(1'h0)] forvar336 = (1'h0);
  reg [(3'h5):(1'h0)] reg335 = (1'h0);
  reg [(5'h17):(1'h0)] forvar331 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg330 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg324 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg321 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg320 = (1'h0);
  reg [(2'h2):(1'h0)] reg319 = (1'h0);
  reg [(5'h13):(1'h0)] reg317 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg315 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg314 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg312 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg310 = (1'h0);
  reg [(5'h14):(1'h0)] reg309 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg307 = (1'h0);
  reg [(4'hb):(1'h0)] forvar306 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg305 = (1'h0);
  reg [(4'h9):(1'h0)] reg304 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar303 = (1'h0);
  reg [(4'he):(1'h0)] forvar302 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg300 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar298 = (1'h0);
  reg [(5'h18):(1'h0)] reg297 = (1'h0);
  reg [(3'h5):(1'h0)] reg296 = (1'h0);
  reg [(5'h13):(1'h0)] reg295 = (1'h0);
  reg [(4'h8):(1'h0)] reg290 = (1'h0);
  reg [(4'h8):(1'h0)] forvar289 = (1'h0);
  reg signed [(5'h15):(1'h0)] forvar287 = (1'h0);
  reg [(4'he):(1'h0)] reg285 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg282 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg279 = (1'h0);
  reg [(3'h4):(1'h0)] reg278 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg277 = (1'h0);
  reg [(5'h10):(1'h0)] reg275 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg274 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar272 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg270 = (1'h0);
  reg [(5'h11):(1'h0)] reg269 = (1'h0);
  reg [(5'h15):(1'h0)] reg267 = (1'h0);
  reg [(3'h4):(1'h0)] forvar266 = (1'h0);
  reg [(4'hf):(1'h0)] reg265 = (1'h0);
  reg [(2'h2):(1'h0)] reg262 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg261 = (1'h0);
  reg [(4'hb):(1'h0)] forvar255 = (1'h0);
  reg [(4'ha):(1'h0)] reg254 = (1'h0);
  reg [(4'hf):(1'h0)] reg253 = (1'h0);
  reg signed [(4'h8):(1'h0)] forvar252 = (1'h0);
  reg [(4'hf):(1'h0)] forvar247 = (1'h0);
  reg [(4'hc):(1'h0)] reg246 = (1'h0);
  reg signed [(4'he):(1'h0)] reg237 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg250 = (1'h0);
  reg [(5'h12):(1'h0)] forvar246 = (1'h0);
  reg [(4'h8):(1'h0)] reg243 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg241 = (1'h0);
  reg [(4'hc):(1'h0)] reg240 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg239 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg238 = (1'h0);
  reg [(3'h4):(1'h0)] forvar237 = (1'h0);
  reg [(5'h10):(1'h0)] reg236 = (1'h0);
  reg [(4'hf):(1'h0)] reg234 = (1'h0);
  reg [(5'h10):(1'h0)] reg229 = (1'h0);
  reg [(5'h10):(1'h0)] forvar223 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg226 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg224 = (1'h0);
  reg [(5'h18):(1'h0)] reg223 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg222 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg218 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg219 = (1'h0);
  reg [(4'h9):(1'h0)] forvar218 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg212 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar203 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg216 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg215 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar212 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg208 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg207 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg206 = (1'h0);
  reg signed [(4'he):(1'h0)] reg202 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg201 = (1'h0);
  assign y = {wire578,
                 wire577,
                 wire575,
                 wire407,
                 wire403,
                 wire402,
                 wire379,
                 wire345,
                 wire323,
                 wire221,
                 wire200,
                 reg203,
                 reg204,
                 reg205,
                 reg209,
                 reg210,
                 reg211,
                 reg213,
                 reg214,
                 reg217,
                 reg220,
                 reg225,
                 reg227,
                 reg228,
                 reg230,
                 reg231,
                 reg232,
                 reg233,
                 reg235,
                 reg242,
                 reg244,
                 reg245,
                 reg247,
                 reg248,
                 reg249,
                 reg251,
                 reg256,
                 reg257,
                 reg258,
                 reg259,
                 reg260,
                 reg263,
                 reg264,
                 reg268,
                 reg271,
                 reg273,
                 reg276,
                 reg280,
                 reg281,
                 reg283,
                 reg284,
                 reg286,
                 reg288,
                 reg291,
                 reg292,
                 reg293,
                 reg294,
                 reg299,
                 reg301,
                 reg308,
                 reg311,
                 reg313,
                 reg316,
                 reg318,
                 reg322,
                 reg325,
                 reg326,
                 reg327,
                 reg328,
                 reg329,
                 reg332,
                 reg333,
                 reg331,
                 reg334,
                 reg337,
                 reg339,
                 reg341,
                 reg336,
                 reg342,
                 reg347,
                 reg348,
                 reg349,
                 reg350,
                 reg351,
                 reg356,
                 reg357,
                 reg359,
                 reg360,
                 reg362,
                 reg363,
                 reg364,
                 reg367,
                 reg369,
                 reg371,
                 reg372,
                 reg373,
                 reg377,
                 reg378,
                 reg382,
                 reg385,
                 reg387,
                 reg384,
                 reg386,
                 reg391,
                 reg395,
                 reg399,
                 reg400,
                 reg404,
                 reg406,
                 reg408,
                 reg409,
                 reg412,
                 reg414,
                 reg419,
                 reg418,
                 reg417,
                 reg416,
                 reg415,
                 reg413,
                 forvar411,
                 forvar410,
                 forvar405,
                 reg401,
                 reg398,
                 forvar397,
                 reg396,
                 reg394,
                 reg393,
                 forvar392,
                 forvar390,
                 reg389,
                 reg388,
                 forvar386,
                 forvar384,
                 reg383,
                 reg381,
                 reg380,
                 forvar376,
                 reg375,
                 reg374,
                 reg370,
                 reg368,
                 reg366,
                 reg365,
                 reg361,
                 reg358,
                 reg355,
                 reg354,
                 reg353,
                 reg352,
                 forvar346,
                 reg344,
                 reg343,
                 reg340,
                 reg338,
                 forvar336,
                 reg335,
                 forvar331,
                 reg330,
                 reg324,
                 reg321,
                 reg320,
                 reg319,
                 reg317,
                 reg315,
                 reg314,
                 reg312,
                 reg310,
                 reg309,
                 reg307,
                 forvar306,
                 reg305,
                 reg304,
                 forvar303,
                 forvar302,
                 reg300,
                 forvar298,
                 reg297,
                 reg296,
                 reg295,
                 reg290,
                 forvar289,
                 forvar287,
                 reg285,
                 reg282,
                 reg279,
                 reg278,
                 reg277,
                 reg275,
                 reg274,
                 forvar272,
                 reg270,
                 reg269,
                 reg267,
                 forvar266,
                 reg265,
                 reg262,
                 reg261,
                 forvar255,
                 reg254,
                 reg253,
                 forvar252,
                 forvar247,
                 reg246,
                 reg237,
                 reg250,
                 forvar246,
                 reg243,
                 reg241,
                 reg240,
                 reg239,
                 reg238,
                 forvar237,
                 reg236,
                 reg234,
                 reg229,
                 forvar223,
                 reg226,
                 reg224,
                 reg223,
                 reg222,
                 reg218,
                 reg219,
                 forvar218,
                 reg212,
                 forvar203,
                 reg216,
                 reg215,
                 forvar212,
                 reg208,
                 reg207,
                 reg206,
                 reg202,
                 reg201,
                 (1'h0)};
  assign wire200 = (~|((~^{$signed(wire199), (!wire199)}) ?
                       wire197[(5'h15):(1'h1)] : wire198[(1'h1):(1'h0)]));
  always
    @(posedge clk) begin
      reg201 = $unsigned($unsigned((~$unsigned(wire196[(1'h0):(1'h0)]))));
      if ($unsigned(($signed(wire197[(3'h4):(2'h2)]) ?
          wire200[(3'h5):(3'h5)] : reg201)))
        begin
          if ($unsigned($unsigned(wire200)))
            begin
              reg202 = $signed($signed($unsigned((&(&wire197)))));
            end
          else
            begin
              reg203 <= (&($signed($signed((wire200 & reg201))) ?
                  reg202[(4'h8):(1'h0)] : wire199[(2'h2):(2'h2)]));
              reg204 <= ({$signed((^wire200)),
                  reg203[(2'h2):(1'h1)]} ~^ {reg201[(2'h3):(1'h1)],
                  (^((reg201 ^~ reg201) <= $unsigned(wire198)))});
            end
          if (reg201)
            begin
              reg205 <= $signed({{(wire199[(1'h1):(1'h0)] && {reg204})}});
              reg206 = $unsigned($signed($unsigned(wire200)));
              reg207 = reg205;
              reg208 = (~|$unsigned(((8'hac) ?
                  $signed((~&wire198)) : ((~|reg203) ^ (!(8'hbf))))));
              reg209 <= (((8'hae) <<< $signed(reg205)) ?
                  (&(&wire199[(2'h2):(1'h1)])) : reg201);
            end
          else
            begin
              reg205 <= $unsigned(wire196[(2'h3):(1'h1)]);
              reg206 = ($signed(reg202[(2'h2):(1'h1)]) - ($signed($unsigned(((8'haf) ?
                  wire199 : (8'ha5)))) ^ $signed(({wire199, reg201} ?
                  $signed(reg205) : wire199[(1'h1):(1'h1)]))));
              reg209 <= (|reg208);
              reg210 <= $unsigned(({(~(^reg209)),
                      $signed((reg208 ? reg204 : reg208))} ?
                  $signed($unsigned((wire196 ?
                      (8'ha4) : reg202))) : (reg203[(2'h2):(2'h2)] ?
                      ($signed(reg206) ?
                          reg204[(3'h5):(2'h3)] : reg207[(3'h7):(3'h5)]) : {(reg201 || wire199)})));
            end
          reg211 <= $unsigned($signed($signed($signed(wire200))));
          for (forvar212 = (1'h0); (forvar212 < (2'h3)); forvar212 = (forvar212 + (1'h1)))
            begin
              reg213 <= (reg210[(4'hb):(3'h7)] * $unsigned(reg205[(1'h1):(1'h1)]));
              reg214 <= (^~($unsigned((((8'ha0) ? reg209 : (8'hb3)) ?
                  (wire196 ? (8'ha6) : wire198) : (reg208 ?
                      forvar212 : (8'hba)))) - (|$unsigned((8'hb7)))));
              reg215 = $unsigned({(((~reg214) - $signed(wire199)) != $signed($signed(wire196)))});
              reg216 = $signed(reg205[(4'hb):(1'h0)]);
              reg217 <= ($signed($unsigned(wire196[(2'h3):(1'h1)])) ?
                  $signed((8'hbd)) : (~^$unsigned(wire196)));
            end
        end
      else
        begin
          reg202 = (8'hb7);
          for (forvar203 = (1'h0); (forvar203 < (1'h1)); forvar203 = (forvar203 + (1'h1)))
            begin
              reg206 = reg216;
              reg207 = reg201[(2'h3):(1'h1)];
              reg209 <= ((reg207[(2'h2):(1'h1)] ~^ $signed(reg213)) ?
                  {(8'ha9),
                      ((!reg206[(1'h1):(1'h0)]) * {wire200[(1'h1):(1'h0)],
                          reg207[(1'h1):(1'h0)]})} : wire199[(1'h1):(1'h1)]);
              reg212 = $unsigned(wire198[(2'h3):(1'h1)]);
              reg213 <= $signed(reg201[(2'h3):(1'h0)]);
            end
        end
      if ((reg202[(4'h8):(4'h8)] >>> $unsigned((($signed(reg216) ?
              $signed(reg208) : reg215) ?
          $unsigned((reg202 ? reg209 : (7'h48))) : (((8'hbf) ?
              wire200 : (8'hb6)) >>> {(7'h49), wire199})))))
        begin
          for (forvar218 = (1'h0); (forvar218 < (1'h1)); forvar218 = (forvar218 + (1'h1)))
            begin
              reg219 = $signed((({$unsigned(reg205)} ?
                  $unsigned((reg207 >= (8'hb9))) : $unsigned($unsigned(reg215))) >= (forvar218 | (reg208[(2'h2):(2'h2)] ?
                  (!(8'ha9)) : $unsigned(wire197)))));
            end
        end
      else
        begin
          reg218 = (^$unsigned(({(reg219 ? wire197 : reg214),
                  $unsigned(reg204)} ?
              {reg205[(2'h2):(1'h1)]} : (~(wire198 >>> forvar218)))));
        end
      reg220 <= reg216;
    end
  assign wire221 = $signed($unsigned({$unsigned((wire196 ?
                           (8'ha6) : reg220))}));
  always
    @(posedge clk) begin
      if ((&reg203))
        begin
          reg222 = (reg211 ?
              ((((reg210 || reg211) ?
                      (+reg211) : $signed(reg214)) >>> $signed({reg217})) ?
                  wire221 : $signed({$signed(reg209)})) : $unsigned(($signed($unsigned(reg204)) ?
                  ($signed(wire200) ?
                      ((8'h9f) || reg203) : {reg220}) : $signed((wire221 ?
                      wire196 : (8'h9f))))));
          reg223 = ((($unsigned({wire221}) ? (|$unsigned(wire221)) : wire221) ?
              (~((reg204 >= wire200) & (wire221 ?
                  reg222 : reg205))) : (~wire199)) >>> $unsigned(wire197));
          if ($unsigned(($unsigned(reg211[(3'h7):(3'h6)]) > $unsigned({$signed(wire199),
              (-wire196)}))))
            begin
              reg224 = wire197;
              reg225 <= {((-(~|{(8'hac)})) >>> reg224), wire197[(4'hc):(4'h9)]};
              reg226 = ($unsigned((($signed(reg209) ?
                  wire199 : $signed(wire221)) << ((reg210 ? wire198 : reg224) ?
                  $unsigned(reg214) : (reg225 ^~ reg213)))) ^ wire197[(1'h0):(1'h0)]);
              reg227 <= (reg204 ~^ $unsigned((reg220 | (8'ha6))));
              reg228 <= (reg209 >= reg210);
            end
          else
            begin
              reg224 = reg203[(2'h2):(1'h1)];
              reg226 = (!($unsigned((+reg226[(5'h14):(5'h12)])) ?
                  (($signed(reg213) >= $signed(reg227)) ?
                      (reg210[(1'h1):(1'h0)] ?
                          (~^wire198) : $signed((7'h46))) : ((wire199 >> reg204) | {reg226})) : ($unsigned($unsigned(reg224)) ?
                      reg227 : wire197)));
            end
        end
      else
        begin
          reg222 = (+($unsigned(reg228) ?
              (wire221[(1'h1):(1'h1)] > reg226) : $signed($unsigned($unsigned(wire198)))));
          for (forvar223 = (1'h0); (forvar223 < (1'h0)); forvar223 = (forvar223 + (1'h1)))
            begin
              reg225 <= {(|(wire200 <<< $unsigned((wire197 ?
                      reg217 : (8'hb6))))),
                  reg220[(2'h2):(1'h1)]};
              reg227 <= forvar223[(2'h2):(1'h1)];
              reg229 = (~^$signed(($signed((reg220 <<< reg209)) & ((~reg204) | $signed(reg209)))));
            end
        end
    end
  always
    @(posedge clk) begin
      if (wire221[(1'h1):(1'h0)])
        begin
          if ((&($signed((^~$unsigned(wire221))) ?
              reg211 : {$signed(wire198[(3'h6):(1'h1)])})))
            begin
              reg230 <= {(8'hb0)};
              reg231 <= (($signed(((reg217 ?
                      reg203 : reg205) ^ wire221[(1'h0):(1'h0)])) >> (8'hb7)) ?
                  (~&(~&$unsigned(reg227[(4'hc):(1'h1)]))) : $signed((({(8'hbb),
                      reg205} ^~ $unsigned(reg205)) != (7'h45))));
            end
          else
            begin
              reg230 <= reg231[(3'h4):(2'h3)];
              reg231 <= (!$signed($signed(wire197[(4'h8):(3'h6)])));
            end
          if (reg211[(3'h5):(2'h2)])
            begin
              reg232 <= {reg231};
              reg233 <= wire198[(3'h6):(1'h1)];
              reg234 = ($signed($unsigned((7'h43))) ?
                  $signed(reg227[(5'h13):(2'h3)]) : {reg210[(4'h9):(3'h6)],
                      (-(wire199[(2'h2):(1'h0)] > reg227[(4'he):(4'he)]))});
              reg235 <= (($unsigned(($unsigned(reg209) ^ $unsigned(reg233))) ?
                      reg213[(3'h5):(1'h1)] : (($signed(reg205) ^~ $signed(reg230)) ?
                          $signed({reg225,
                              wire221}) : (reg227 - $unsigned(reg225)))) ?
                  (&$unsigned(($unsigned(reg234) > reg203))) : wire221);
            end
          else
            begin
              reg234 = reg205[(4'h9):(3'h6)];
              reg236 = ($signed(reg211[(4'hb):(3'h7)]) ?
                  reg227 : $signed(wire199[(1'h0):(1'h0)]));
            end
        end
      else
        begin
          reg234 = ($unsigned(wire221) ?
              (reg228[(2'h2):(1'h0)] ^~ wire221[(1'h0):(1'h0)]) : $signed((((~&reg217) ?
                      reg231 : (reg217 == wire196)) ?
                  reg230[(4'hb):(4'h8)] : $signed({reg233, reg220}))));
          reg236 = wire197;
        end
      if ((reg235 || $signed($unsigned((~^$signed(reg220))))))
        begin
          for (forvar237 = (1'h0); (forvar237 < (2'h2)); forvar237 = (forvar237 + (1'h1)))
            begin
              reg238 = $unsigned($signed(((~reg214[(5'h11):(5'h11)]) == reg210)));
            end
          reg239 = {($signed((~&$signed((8'hb1)))) ?
                  reg220[(2'h2):(2'h2)] : $signed(reg214))};
          if (reg205[(3'h6):(3'h4)])
            begin
              reg240 = (((reg239[(1'h0):(1'h0)] > (8'ha0)) ?
                  wire221[(1'h1):(1'h0)] : $signed(reg209[(3'h5):(2'h3)])) < reg214[(4'hc):(3'h5)]);
              reg241 = $signed(reg233[(4'hb):(1'h1)]);
              reg242 <= ($signed($signed((reg236 >> (reg225 ^~ (8'hbd))))) ?
                  {$signed(($unsigned(reg240) ? {wire221} : (^reg239))),
                      {$signed((8'ha4)),
                          reg217[(3'h4):(2'h3)]}} : (^~(reg238 <= reg233[(3'h5):(1'h1)])));
              reg243 = $signed(reg210[(3'h7):(3'h6)]);
              reg244 <= (reg214[(1'h0):(1'h0)] >>> {$unsigned($unsigned(((8'hac) & reg210))),
                  $signed((~$signed(reg240)))});
            end
          else
            begin
              reg242 <= $signed(reg213);
              reg243 = (8'hae);
              reg244 <= $signed((8'haa));
              reg245 <= $signed((7'h47));
            end
          for (forvar246 = (1'h0); (forvar246 < (1'h0)); forvar246 = (forvar246 + (1'h1)))
            begin
              reg247 <= (!(($unsigned({reg234,
                  reg231}) <= (^~(+wire198))) >> $unsigned((-(8'had)))));
              reg248 <= (-reg236);
              reg249 <= $unsigned($unsigned((+reg248[(5'h10):(4'hb)])));
            end
          reg250 = $unsigned({($unsigned(wire199[(2'h2):(1'h0)]) ?
                  reg244 : wire221)});
        end
      else
        begin
          reg237 = $unsigned({wire196, (!$signed($unsigned(wire197)))});
          if (reg205)
            begin
              reg238 = wire197[(4'hf):(2'h3)];
              reg239 = reg209[(1'h1):(1'h1)];
            end
          else
            begin
              reg238 = reg249;
              reg239 = ($unsigned((~^(reg210 * reg217[(2'h3):(1'h0)]))) ?
                  $unsigned({((reg236 <= reg235) ?
                          {reg203} : (~reg205))}) : reg211[(3'h6):(3'h5)]);
              reg242 <= (reg247[(4'ha):(1'h1)] ?
                  reg238[(3'h6):(1'h0)] : $signed((8'haa)));
              reg244 <= reg244[(5'h11):(1'h1)];
              reg245 <= (~^(({{reg233, wire197}, $signed(reg205)} ?
                  reg234 : reg238[(3'h4):(1'h1)]) > (~{$signed((8'hab))})));
            end
          reg246 = $signed($signed($signed($unsigned((reg242 <<< reg247)))));
          for (forvar247 = (1'h0); (forvar247 < (2'h3)); forvar247 = (forvar247 + (1'h1)))
            begin
              reg248 <= (reg246[(4'ha):(2'h3)] ?
                  reg245[(3'h6):(2'h2)] : $unsigned(((reg240[(4'h8):(2'h3)] ?
                          (reg211 ? reg248 : reg205) : $signed(reg228)) ?
                      $signed({reg244}) : reg248[(4'hb):(2'h3)])));
              reg250 = $unsigned(reg204[(2'h2):(1'h0)]);
            end
        end
      reg251 <= $signed(((~&{(reg246 >>> reg234)}) ^ (reg237 ?
          $signed((|(7'h42))) : (8'haf))));
      for (forvar252 = (1'h0); (forvar252 < (2'h3)); forvar252 = (forvar252 + (1'h1)))
        begin
          reg253 = $signed((reg228[(4'ha):(3'h7)] >> {(!(^forvar247)),
              ((^reg242) ? reg233 : {reg247, reg237})}));
          reg254 = (^~{(-{(reg241 ? reg211 : reg203)}),
              wire197[(4'ha):(3'h7)]});
          for (forvar255 = (1'h0); (forvar255 < (2'h2)); forvar255 = (forvar255 + (1'h1)))
            begin
              reg256 <= ((&{(^~reg242)}) && $signed((reg245[(2'h2):(2'h2)] + (!$signed(reg238)))));
              reg257 <= reg220[(2'h2):(1'h1)];
              reg258 <= $signed(((8'hb0) ?
                  (&{(forvar255 >> reg227)}) : ($signed((^~(7'h42))) - $unsigned(reg250))));
              reg259 <= wire199;
              reg260 <= reg238[(2'h2):(1'h1)];
            end
          if ((reg241[(3'h5):(3'h5)] ?
              forvar246[(4'hc):(4'ha)] : (((~|(^~reg253)) ?
                      $unsigned((~&(8'hb7))) : ($unsigned(reg211) ~^ $unsigned(reg250))) ?
                  reg256[(4'hb):(2'h3)] : $signed(((reg244 ?
                      reg257 : (8'h9e)) <= (forvar252 && reg228))))))
            begin
              reg261 = reg240[(1'h1):(1'h1)];
              reg262 = (~^((forvar252[(1'h1):(1'h1)] + $signed($signed(reg230))) == {$unsigned((reg203 ?
                      reg205 : reg225)),
                  reg214}));
              reg263 <= $unsigned($signed($unsigned(((|reg256) << $signed(reg214)))));
              reg264 <= (+{(reg263 << $signed($unsigned((8'hb4))))});
              reg265 = ((wire196[(3'h5):(2'h2)] | (!(reg211[(4'hf):(3'h6)] ?
                      ((8'hb6) ? reg243 : reg260) : (reg231 ?
                          (8'hb7) : reg246)))) ?
                  $signed(($unsigned($signed(reg251)) >>> $signed($signed(reg242)))) : (-$unsigned(reg239[(4'hb):(3'h7)])));
            end
          else
            begin
              reg261 = $unsigned(reg231[(1'h1):(1'h0)]);
              reg263 <= reg261[(4'h8):(3'h5)];
            end
          for (forvar266 = (1'h0); (forvar266 < (3'h4)); forvar266 = (forvar266 + (1'h1)))
            begin
              reg267 = $signed(reg262);
              reg268 <= (|$unsigned($signed((~^$unsigned(reg267)))));
              reg269 = $signed(($signed(reg243) >>> (reg243 == $unsigned(reg241))));
              reg270 = $signed($unsigned($unsigned(($signed(reg227) ?
                  reg210 : $signed(wire221)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg271 <= reg263;
      for (forvar272 = (1'h0); (forvar272 < (3'h4)); forvar272 = (forvar272 + (1'h1)))
        begin
          reg273 <= wire198;
          reg274 = ((-($signed(reg263[(1'h0):(1'h0)]) >> ($signed((8'h9d)) ?
                  (&reg273) : {reg211}))) ?
              $signed((~&(7'h4a))) : ($unsigned(((reg256 == reg256) | $unsigned(reg249))) > $signed(reg203)));
          reg275 = reg263[(1'h1):(1'h0)];
        end
      if ((((((~&reg233) ~^ $signed(forvar272)) != {((8'h9c) ?
                  reg225 : reg268)}) - (~|reg227[(5'h15):(5'h15)])) ?
          $signed($signed($unsigned((wire200 ?
              (8'hb6) : reg203)))) : $signed($signed($signed(reg257)))))
        begin
          reg276 <= $signed(wire198);
          if (reg209[(4'hf):(4'hb)])
            begin
              reg277 = {$signed(reg211)};
              reg278 = ($unsigned((reg232 ?
                  wire198[(2'h2):(1'h0)] : wire200)) & $unsigned(((~^(reg276 & reg273)) ?
                  $unsigned((!(8'hb5))) : reg231)));
              reg279 = reg251;
            end
          else
            begin
              reg277 = $signed(reg231[(1'h1):(1'h0)]);
              reg278 = ($signed($unsigned((^(~|reg244)))) * reg209);
              reg280 <= (({$signed((wire197 ? (8'hac) : reg210)),
                  ((~|reg256) ?
                      reg268 : $signed(reg209))} ^~ (~&(~reg245[(1'h1):(1'h0)]))) != $signed({($signed(reg205) >>> (|reg244)),
                  forvar272[(1'h1):(1'h0)]}));
            end
          if (($unsigned($signed(reg245)) ?
              $unsigned(wire200) : ($unsigned(reg230[(3'h6):(1'h1)]) ?
                  reg263 : $signed({(reg211 == reg244), (~|wire198)}))))
            begin
              reg281 <= (reg268[(4'hd):(4'h8)] >> $unsigned((!((reg230 ?
                      reg225 : (8'hba)) ?
                  $signed(reg280) : $unsigned(reg232)))));
              reg282 = (reg204[(1'h0):(1'h0)] ?
                  $signed({(^((8'ha5) ?
                          reg264 : reg259))}) : $signed($unsigned(reg275)));
              reg283 <= (~(($unsigned((reg259 == (8'hac))) <<< reg251[(3'h4):(1'h0)]) ?
                  $unsigned($signed((^reg230))) : $signed($signed({(8'hb1)}))));
              reg284 <= (reg203[(2'h2):(1'h0)] >= wire200[(2'h3):(2'h3)]);
            end
          else
            begin
              reg281 <= (((~&reg231[(3'h4):(1'h0)]) ?
                      $signed($signed((reg227 | (8'hb9)))) : $signed((|{reg228}))) ?
                  (~^$signed(((reg258 | (8'ha9)) * reg231))) : ((($unsigned((8'ha6)) ?
                          (reg233 >= reg228) : {reg263}) + ({reg225, reg256} ?
                          reg217 : (reg260 ? (8'h9c) : wire198))) ?
                      reg249 : $unsigned(reg268[(3'h7):(3'h6)])));
              reg283 <= reg231[(4'h8):(1'h1)];
              reg285 = reg227;
            end
          reg286 <= {((reg247[(3'h4):(2'h3)] <<< reg233[(5'h14):(4'hb)]) ?
                  $signed((|reg264[(2'h2):(1'h1)])) : $signed($unsigned((reg260 << reg273))))};
        end
      else
        begin
          reg277 = reg275;
        end
      for (forvar287 = (1'h0); (forvar287 < (3'h4)); forvar287 = (forvar287 + (1'h1)))
        begin
          reg288 <= (^~((reg258[(2'h2):(1'h1)] ?
              ((8'hbd) || wire199[(2'h2):(1'h1)]) : (+reg245)) || (~|(reg282[(4'h8):(1'h0)] <<< reg205[(4'ha):(3'h6)]))));
          for (forvar289 = (1'h0); (forvar289 < (1'h1)); forvar289 = (forvar289 + (1'h1)))
            begin
              reg290 = (reg271 ^ (({$unsigned(reg244)} ?
                      (reg214[(4'hb):(3'h7)] ?
                          reg277[(5'h14):(4'hb)] : reg217[(1'h1):(1'h0)]) : $signed($unsigned(reg280))) ?
                  (((!forvar272) ?
                      {reg288,
                          reg247} : (reg257 ^ reg273)) && reg249) : reg231));
              reg291 <= ((8'hac) ?
                  $signed((((reg259 ? reg214 : reg271) == (reg242 ?
                      wire197 : reg247)) | (reg247[(4'h9):(3'h6)] > $signed(reg281)))) : ($unsigned($unsigned($signed((8'ha6)))) <= $signed({{wire197,
                          reg209}})));
              reg292 <= ((~^($signed($signed(reg245)) != reg227)) ?
                  wire198[(4'h8):(3'h4)] : (~reg257[(2'h3):(2'h2)]));
            end
          if (($unsigned(($signed((~&reg280)) < $signed((reg263 ?
                  reg249 : reg209)))) ?
              {{$unsigned($unsigned(reg257))},
                  reg280} : ($signed((^~$unsigned(reg292))) ?
                  $signed(reg276) : {(~reg292)})))
            begin
              reg293 <= (~|{$signed({$signed(reg217)})});
              reg294 <= $signed(reg257);
            end
          else
            begin
              reg295 = (^$signed(((~((8'hac) ?
                  reg263 : reg256)) - $unsigned($unsigned(wire199)))));
              reg296 = {(~^reg225)};
              reg297 = {$unsigned(($signed(wire200) == reg284)),
                  reg232[(2'h3):(2'h2)]};
            end
        end
      for (forvar298 = (1'h0); (forvar298 < (2'h2)); forvar298 = (forvar298 + (1'h1)))
        begin
          reg299 <= $unsigned(reg251[(1'h1):(1'h0)]);
          reg300 = $unsigned(reg281[(5'h16):(5'h13)]);
          reg301 <= {reg235};
        end
    end
  always
    @(posedge clk) begin
      for (forvar302 = (1'h0); (forvar302 < (2'h3)); forvar302 = (forvar302 + (1'h1)))
        begin
          for (forvar303 = (1'h0); (forvar303 < (2'h3)); forvar303 = (forvar303 + (1'h1)))
            begin
              reg304 = reg280;
              reg305 = {{reg299[(3'h6):(1'h0)],
                      $signed(({reg284, reg204} ?
                          reg258[(3'h4):(2'h2)] : reg230))}};
            end
          for (forvar306 = (1'h0); (forvar306 < (2'h2)); forvar306 = (forvar306 + (1'h1)))
            begin
              reg307 = reg263;
              reg308 <= $signed(((+{$signed(reg227),
                  $signed(reg242)}) >>> reg268[(2'h3):(1'h0)]));
            end
        end
      if ($unsigned(wire198))
        begin
          if ((-reg305))
            begin
              reg309 = (~&(reg260[(4'hc):(2'h2)] || forvar306[(1'h1):(1'h1)]));
              reg310 = ($unsigned({(reg283 - (+reg301))}) ?
                  $unsigned(((-$signed(reg245)) ^ (reg228[(4'h9):(1'h0)] ?
                      $unsigned(reg308) : ((7'h45) ?
                          (8'hb5) : wire197)))) : $unsigned($signed($unsigned((&(8'ha6))))));
              reg311 <= ((reg307[(3'h7):(3'h4)] ?
                  reg209[(3'h5):(1'h0)] : (reg310[(3'h7):(3'h5)] >> $unsigned((wire199 ^ reg310)))) ^~ $signed($unsigned($unsigned((reg204 ?
                  reg291 : reg213)))));
              reg312 = (reg245[(4'h8):(2'h2)] * $signed(reg291));
              reg313 <= (-($signed((&$signed(reg220))) & $unsigned(((reg220 >>> reg231) + reg284[(4'ha):(4'h8)]))));
            end
          else
            begin
              reg309 = (~forvar302);
              reg310 = reg311[(3'h7):(1'h1)];
              reg311 <= (8'ha6);
              reg312 = (($unsigned($signed((reg304 == (8'hbe)))) && reg313[(4'h8):(1'h0)]) ?
                  ($signed(reg308[(3'h4):(2'h3)]) >> reg312[(4'h8):(2'h2)]) : ((((reg211 * wire200) > (8'haa)) ?
                      wire200[(3'h4):(2'h3)] : (reg242[(4'hd):(2'h2)] ?
                          $unsigned(reg259) : (reg227 ?
                              reg313 : reg220))) < $signed(($signed(reg312) ?
                      $unsigned((8'hba)) : (reg245 ? reg258 : reg301)))));
            end
          reg314 = (reg213 >> ((^~$unsigned(reg233)) ~^ (^(wire198 || reg299[(2'h2):(1'h1)]))));
        end
      else
        begin
          reg311 <= (|(reg256[(5'h11):(3'h6)] ?
              (reg258[(2'h3):(2'h2)] ?
                  $unsigned(((8'hb1) | (8'ha0))) : $unsigned((~reg299))) : ($unsigned((wire199 && reg292)) ?
                  ((reg311 ?
                      forvar302 : reg293) || $signed((7'h4a))) : ({(7'h48)} + forvar302))));
          reg313 <= $signed(($signed(reg309) ?
              $signed(reg257) : $signed((~(~|(8'hbb))))));
          reg314 = {wire198, $unsigned((~&reg263[(1'h0):(1'h0)]))};
          reg315 = $signed(($signed($signed($unsigned(reg235))) * $unsigned(reg225[(1'h1):(1'h1)])));
          if ($signed((~^$signed((^(reg307 ? reg249 : reg309))))))
            begin
              reg316 <= $unsigned($signed((|reg209[(2'h2):(1'h0)])));
              reg317 = $unsigned(reg235[(5'h10):(4'hb)]);
              reg318 <= (8'ha3);
              reg319 = {wire198[(1'h0):(1'h0)], reg235};
              reg320 = (8'hb1);
            end
          else
            begin
              reg316 <= reg304[(3'h5):(2'h3)];
            end
        end
      reg321 = $unsigned($signed((~&$signed($unsigned(reg273)))));
      reg322 <= $signed(wire197);
    end
  assign wire323 = reg217[(5'h12):(5'h12)];
  always
    @(posedge clk) begin
      if (reg308[(2'h3):(1'h1)])
        begin
          reg324 = $signed(($unsigned(wire197) ?
              $signed(((reg322 >>> reg227) >= ((8'hbe) ?
                  reg276 : reg286))) : ({(~&reg273), (~&reg293)} <= (7'h40))));
          if ($unsigned(($signed(({(7'h44)} | ((8'ha6) ?
              (8'ha7) : reg245))) > (~^reg301[(1'h1):(1'h1)]))))
            begin
              reg325 <= {(~(8'hb2)), $unsigned($unsigned($unsigned(reg260)))};
              reg326 <= ({$signed(($unsigned(reg280) ?
                          (reg220 ^ reg251) : reg217)),
                      $unsigned($unsigned($signed(reg235)))} ?
                  reg227[(3'h4):(2'h2)] : (reg308[(2'h2):(1'h1)] ?
                      $unsigned(reg263) : ($unsigned($signed(reg209)) << $unsigned(((7'h40) ?
                          reg259 : reg311)))));
              reg327 <= ($signed(($signed(reg244) ?
                  (8'hbf) : reg210)) <= $unsigned((|(8'hb8))));
              reg328 <= reg217;
              reg329 <= $signed($unsigned(($signed($signed(wire200)) ~^ $signed(reg245[(1'h1):(1'h0)]))));
            end
          else
            begin
              reg330 = ($signed((&{(reg327 <= reg231)})) ?
                  ($signed((~&(^~reg248))) > $signed(reg213)) : (((^$unsigned(reg271)) <= reg204) ?
                      $signed(reg251) : (+($signed(reg245) ^~ $signed(reg258)))));
            end
          for (forvar331 = (1'h0); (forvar331 < (1'h1)); forvar331 = (forvar331 + (1'h1)))
            begin
              reg332 <= {((((reg268 + reg232) << (reg271 ?
                      reg225 : (8'ha7))) ^ reg268[(4'h9):(4'h8)]) << ((^(8'hbb)) ?
                      $unsigned(reg268) : reg271)),
                  $unsigned($signed((+$signed((8'hbf)))))};
              reg333 <= ($signed((&(reg276[(4'h9):(4'h9)] ?
                  $signed((8'hbe)) : (&reg242)))) != reg204);
            end
        end
      else
        begin
          reg325 <= reg293;
          reg326 <= ($unsigned($signed($signed(wire200))) <= $signed(((~&$unsigned(reg276)) >> $unsigned(reg324))));
          reg330 = {reg326};
          reg331 <= $unsigned(reg264);
        end
      reg334 <= reg271[(5'h13):(2'h3)];
    end
  always
    @(posedge clk) begin
      reg335 = $signed((($signed($signed(wire199)) ?
              $signed($unsigned(reg284)) : $signed($unsigned(reg248))) ?
          (-((wire198 && (8'ha2)) ?
              reg268[(3'h5):(2'h2)] : (~&reg248))) : $signed($unsigned(reg205))));
      if ($unsigned((~^$signed($signed(reg326[(1'h1):(1'h0)])))))
        begin
          for (forvar336 = (1'h0); (forvar336 < (3'h4)); forvar336 = (forvar336 + (1'h1)))
            begin
              reg337 <= reg247[(2'h3):(1'h0)];
              reg338 = $signed(reg264[(3'h5):(2'h2)]);
              reg339 <= $signed(reg288);
              reg340 = $unsigned(reg280);
              reg341 <= ((^$signed($signed((reg204 && reg256)))) ?
                  $unsigned((&$signed((reg209 == reg204)))) : reg326[(4'h8):(3'h4)]);
            end
        end
      else
        begin
          reg336 <= ($unsigned($unsigned((!$unsigned(reg220)))) < $signed(reg220[(4'hc):(3'h5)]));
          reg338 = $unsigned($unsigned((((~^reg288) | $unsigned(reg281)) ?
              ((~reg245) <<< (!reg228)) : $signed(reg329[(1'h0):(1'h0)]))));
        end
      reg342 <= $unsigned((~^{$signed((reg313 ? (8'hac) : reg244))}));
      reg343 = ($signed($unsigned(((reg313 <= reg342) ?
          $unsigned((8'h9e)) : (7'h41)))) <<< (|($unsigned((!wire221)) ?
          (~((7'h44) ? reg284 : reg233)) : wire221[(1'h0):(1'h0)])));
    end
  always
    @(posedge clk) begin
      reg344 = reg263;
    end
  assign wire345 = (^({(~&wire197[(1'h1):(1'h0)]),
                           ((reg264 ? reg264 : reg225) ?
                               reg284 : (reg227 <= reg268))} ?
                       reg325 : reg230[(3'h7):(3'h4)]));
  always
    @(posedge clk) begin
      if (reg337)
        begin
          for (forvar346 = (1'h0); (forvar346 < (3'h4)); forvar346 = (forvar346 + (1'h1)))
            begin
              reg347 <= $signed(reg301);
              reg348 <= ((!{$signed((reg276 + reg329)),
                      ($unsigned(reg333) ? $signed(reg256) : reg210)}) ?
                  (reg258[(3'h4):(3'h4)] ?
                      (($signed(reg292) * $signed(reg264)) != ((reg210 != reg248) - reg248)) : reg263[(2'h2):(1'h0)]) : ({$unsigned(((7'h45) ^ reg337)),
                          (|(reg220 || wire199))} ?
                      wire323 : reg203));
              reg349 <= (~|wire196);
              reg350 <= (+($signed((~|(reg337 & reg334))) ?
                  reg227[(1'h0):(1'h0)] : (|wire221[(1'h0):(1'h0)])));
            end
          reg351 <= reg350[(5'h10):(2'h2)];
        end
      else
        begin
          for (forvar346 = (1'h0); (forvar346 < (1'h1)); forvar346 = (forvar346 + (1'h1)))
            begin
              reg352 = ((reg244[(3'h4):(1'h1)] ^ (((reg211 == reg248) + {reg256,
                  reg339}) ~^ reg341)) & ($signed(({reg205,
                  reg316} < $unsigned(reg205))) >> {reg342[(4'h9):(3'h5)],
                  ({reg210, reg350} ? reg291 : $signed(reg256))}));
              reg353 = reg231;
              reg354 = ($unsigned((~|(reg288 ?
                  reg322 : (!reg256)))) << $signed($signed($unsigned(reg334))));
            end
          if ($unsigned(reg217[(5'h15):(3'h7)]))
            begin
              reg355 = reg311;
            end
          else
            begin
              reg356 <= {$unsigned((~|$unsigned(reg351))), $unsigned({reg291})};
              reg357 <= reg308[(2'h2):(2'h2)];
            end
        end
      reg358 = reg281;
      reg359 <= $unsigned((reg283[(1'h1):(1'h1)] - ((~|reg271) >> ($signed(reg311) & (reg288 < reg316)))));
      if (((+({(+reg235),
          $signed((8'hac))} <<< $signed($signed(reg280)))) < reg228))
        begin
          if ((~^reg313[(4'h9):(3'h6)]))
            begin
              reg360 <= $signed(wire200);
              reg361 = (8'h9f);
              reg362 <= $signed(reg329);
              reg363 <= $unsigned(($unsigned(({reg347, reg228} > reg354)) ?
                  (-(~^reg331)) : (&((reg316 ? reg301 : wire221) ?
                      $signed(reg358) : $unsigned(reg350)))));
              reg364 <= (-reg256);
            end
          else
            begin
              reg361 = (~((reg359 ?
                      (|$unsigned(wire198)) : (~&(reg203 ? (7'h4a) : reg245))) ?
                  (reg293 ~^ $unsigned((!reg313))) : (((reg349 ?
                          reg337 : reg334) ?
                      (reg220 ?
                          reg358 : reg248) : $unsigned((8'hab))) & ((8'hb3) ^ (reg325 | (8'ha9))))));
              reg365 = (8'hb3);
              reg366 = reg362;
            end
          reg367 <= reg359[(3'h6):(3'h4)];
          if ((&{reg284[(4'ha):(3'h5)], reg325[(3'h5):(2'h3)]}))
            begin
              reg368 = reg367;
              reg369 <= wire200[(3'h7):(3'h6)];
              reg370 = $unsigned($signed((8'hae)));
              reg371 <= (reg362[(1'h1):(1'h1)] ?
                  (reg370[(3'h6):(3'h4)] + ((reg286 ?
                          $unsigned(reg245) : (+reg331)) ?
                      ({reg204,
                          reg281} && $signed(wire200)) : ($signed(reg242) + (~reg291)))) : ($signed($unsigned((reg363 || reg288))) ?
                      {($signed(reg334) ^ reg342[(4'hf):(3'h7)]),
                          (~|reg367[(4'h8):(3'h4)])} : wire345[(3'h7):(3'h7)]));
            end
          else
            begin
              reg368 = reg318;
              reg370 = $signed((reg291[(4'hb):(3'h4)] & reg337));
              reg371 <= ($unsigned(reg364[(4'hc):(2'h3)]) ?
                  (($signed(reg354[(1'h1):(1'h0)]) >= {(&reg328)}) ?
                      (reg329[(1'h0):(1'h0)] << (&{reg233})) : $signed((&reg263[(1'h0):(1'h0)]))) : (+$unsigned(({reg217,
                      reg341} != reg301[(2'h3):(2'h2)]))));
              reg372 <= reg326[(3'h5):(2'h2)];
              reg373 <= (+(reg355 ?
                  reg258[(3'h4):(1'h1)] : reg293[(3'h6):(3'h4)]));
            end
          reg374 = ((~&(reg233 ^ (-reg326[(4'h9):(3'h4)]))) ?
              {reg257[(5'h14):(4'hf)]} : (($unsigned((reg231 ^~ reg231)) * $unsigned($unsigned(reg284))) < reg271[(2'h3):(2'h2)]));
          reg375 = (reg280[(2'h2):(1'h1)] & reg355);
        end
      else
        begin
          if ((~&(&((reg281[(4'hd):(2'h3)] ?
              (8'ha5) : $unsigned(reg276)) && reg271[(4'he):(3'h5)]))))
            begin
              reg361 = $signed(reg231);
            end
          else
            begin
              reg361 = (~^(($signed($unsigned((8'hb1))) * (!(reg329 ?
                      reg363 : reg213))) ?
                  $signed(reg251) : $signed($signed(reg284))));
              reg362 <= (reg374[(5'h11):(4'h8)] ? (!(~|(8'ha1))) : reg359);
              reg365 = (reg260 ?
                  (~^(!{(&(8'hbf)), (!reg375)})) : {reg284,
                      $unsigned($unsigned(reg308[(2'h2):(2'h2)]))});
              reg367 <= ((~^$signed($unsigned({reg351}))) ?
                  $signed(reg249[(2'h3):(1'h1)]) : (&reg359[(3'h4):(3'h4)]));
            end
        end
      for (forvar376 = (1'h0); (forvar376 < (2'h2)); forvar376 = (forvar376 + (1'h1)))
        begin
          reg377 <= $signed(reg244[(3'h6):(2'h3)]);
          reg378 <= (|(reg375[(4'h8):(3'h5)] ~^ reg366));
        end
    end
  assign wire379 = (reg286[(2'h3):(2'h2)] ~^ ((&reg213) ?
                       reg356 : (+($signed((7'h46)) ?
                           {reg205, reg233} : $signed((8'haa))))));
  always
    @(posedge clk) begin
      reg380 = $signed($signed($unsigned(reg230)));
      if ({reg313[(3'h7):(1'h1)], ((!$signed((-reg373))) ^~ wire379)})
        begin
          reg381 = (((8'ha8) ? (~|$unsigned((-reg204))) : (&reg377)) ?
              wire323[(3'h6):(3'h5)] : $signed((reg225 ?
                  {(&reg203)} : ((reg248 ? wire221 : reg230) << (^~reg350)))));
          if ({$unsigned($signed(((reg334 == reg380) ?
                  (reg318 < reg247) : reg233)))})
            begin
              reg382 <= ($signed({reg232[(3'h7):(3'h5)]}) ~^ $signed((~&reg283)));
            end
          else
            begin
              reg383 = $unsigned((&reg292[(4'h8):(3'h7)]));
            end
          for (forvar384 = (1'h0); (forvar384 < (1'h1)); forvar384 = (forvar384 + (1'h1)))
            begin
              reg385 <= (~$unsigned((~reg329[(1'h1):(1'h1)])));
            end
          for (forvar386 = (1'h0); (forvar386 < (1'h0)); forvar386 = (forvar386 + (1'h1)))
            begin
              reg387 <= reg280;
              reg388 = ((($signed({reg359, (8'hb3)}) ?
                      {(wire345 & (8'hb0)),
                          wire323} : $unsigned($unsigned(reg256))) < $signed($unsigned((reg360 ^ reg334)))) ?
                  reg356 : ((reg209[(4'hb):(4'h9)] ?
                      {{reg351},
                          reg260[(4'ha):(3'h4)]} : (^~(~|reg294))) ^~ (+{{reg329,
                          reg337},
                      reg371})));
            end
          reg389 = ((~&(((!reg316) + reg342) == wire221[(1'h1):(1'h1)])) ?
              {wire323, reg362[(2'h2):(1'h0)]} : reg283[(4'ha):(2'h2)]);
        end
      else
        begin
          if (reg214[(4'he):(2'h2)])
            begin
              reg382 <= reg299;
            end
          else
            begin
              reg382 <= reg291;
              reg384 <= ((-wire196) ? reg388[(5'h16):(2'h2)] : reg292);
              reg385 <= ($unsigned(reg204[(3'h6):(2'h2)]) ?
                  reg230 : (!{reg214, reg327}));
              reg386 <= ((reg385[(3'h5):(3'h5)] ?
                      $unsigned((|{reg349})) : ({(8'haf), (~reg235)} ?
                          reg339 : (|reg384[(3'h6):(3'h4)]))) ?
                  reg389[(4'h9):(3'h6)] : reg327);
            end
          reg388 = reg225[(3'h5):(3'h5)];
          reg389 = reg264;
          for (forvar390 = (1'h0); (forvar390 < (1'h1)); forvar390 = (forvar390 + (1'h1)))
            begin
              reg391 <= ((~^reg332[(2'h2):(1'h0)]) ^~ reg257[(5'h10):(2'h3)]);
            end
          for (forvar392 = (1'h0); (forvar392 < (1'h0)); forvar392 = (forvar392 + (1'h1)))
            begin
              reg393 = (((((reg214 ? reg276 : reg308) ^~ (reg339 ?
                  wire200 : reg367)) | wire379[(1'h1):(1'h1)]) >> $unsigned($unsigned($unsigned((7'h41))))) >>> reg227[(3'h7):(3'h4)]);
              reg394 = $unsigned((|reg213));
              reg395 <= reg256;
            end
        end
      reg396 = reg225[(1'h0):(1'h0)];
      for (forvar397 = (1'h0); (forvar397 < (1'h1)); forvar397 = (forvar397 + (1'h1)))
        begin
          if ((7'h40))
            begin
              reg398 = $signed({reg256[(4'h9):(3'h6)], reg211[(3'h7):(2'h3)]});
            end
          else
            begin
              reg399 <= ($unsigned(reg291) ?
                  ((!$unsigned($unsigned(reg318))) ?
                      ((|(reg294 ~^ wire323)) ?
                          reg387 : reg247) : $unsigned($signed((reg339 ?
                          reg331 : (8'hb9))))) : $signed(reg301[(3'h4):(1'h1)]));
            end
          reg400 <= reg299[(3'h5):(1'h1)];
        end
      reg401 = $unsigned((-reg371));
    end
  assign wire402 = (8'hb9);
  assign wire403 = $signed(($signed($signed((~&wire379))) << (reg399 >> {(~|wire200),
                       reg316[(3'h5):(2'h2)]})));
  always
    @(posedge clk) begin
      reg404 <= ($unsigned((&reg286)) ? (!reg281[(5'h15):(3'h7)]) : reg233);
      for (forvar405 = (1'h0); (forvar405 < (2'h2)); forvar405 = (forvar405 + (1'h1)))
        begin
          reg406 <= $signed($unsigned(wire197));
        end
    end
  assign wire407 = reg382[(1'h0):(1'h0)];
  always
    @(posedge clk) begin
      reg408 <= ($unsigned({$signed($signed((8'hb9))),
          $unsigned((reg301 ?
              reg203 : reg230))}) <<< ((~|(&(-(8'hae)))) > ((|(-reg231)) ?
          reg322[(4'hf):(4'h8)] : $unsigned($unsigned(wire200)))));
      reg409 <= $unsigned((|(($unsigned(reg333) ?
          $signed(wire197) : (~&wire221)) > $signed(reg336))));
    end
  always
    @(posedge clk) begin
      for (forvar410 = (1'h0); (forvar410 < (2'h3)); forvar410 = (forvar410 + (1'h1)))
        begin
          for (forvar411 = (1'h0); (forvar411 < (3'h4)); forvar411 = (forvar411 + (1'h1)))
            begin
              reg412 <= wire197;
            end
          reg413 = reg259[(2'h2):(1'h1)];
          if ((-reg247[(3'h7):(1'h1)]))
            begin
              reg414 <= ($unsigned((reg232 ?
                      reg326[(4'h8):(3'h6)] : reg336[(1'h0):(1'h0)])) ?
                  $signed((reg413[(1'h0):(1'h0)] + reg362[(1'h0):(1'h0)])) : $unsigned($unsigned(reg349[(2'h2):(2'h2)])));
            end
          else
            begin
              reg414 <= $signed($signed((((^~reg332) ?
                  {reg367,
                      (8'ha6)} : $unsigned(reg414)) < wire200[(1'h1):(1'h0)])));
              reg415 = reg331[(5'h14):(4'hb)];
              reg416 = $signed(($signed(((wire323 ?
                  reg313 : reg203) && wire198)) & $signed((~|(~^reg286)))));
              reg417 = $signed($unsigned(reg228));
            end
          reg418 = $signed($signed(($unsigned(reg247[(4'ha):(3'h7)]) != ((&reg280) == reg336))));
          reg419 = reg357;
        end
    end
  module420 #() modinst576 (.wire425(reg316), .wire421(reg378), .clk(clk), .wire424(reg384), .y(wire575), .wire422(reg359), .wire423(reg227));
  assign wire577 = (~|($unsigned(((reg399 & reg414) ?
                       $signed(reg339) : reg372[(3'h5):(3'h5)])) ~^ (~^$unsigned((reg334 ^~ reg362)))));
  assign wire578 = $signed($unsigned(reg227));
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module420
#(parameter param574 = (({(((7'h40) + (8'hb4)) < ((7'h41) ? (8'haa) : (7'h42)))} * {((~^(8'ha1)) << ((7'h4a) ^~ (7'h41)))}) ? {(~(((8'haa) ~^ (7'h49)) ? (~|(8'h9d)) : ((8'ha8) & (8'hb0)))), ({((7'h45) ? (8'hac) : (8'ha0)), (-(8'had))} | (^~((8'h9e) ? (8'ha6) : (7'h44))))} : ((+((!(8'hb8)) ? ((8'hb2) ~^ (7'h4a)) : (+(8'ha7)))) ? {(((8'hbd) ? (8'ha0) : (8'ha4)) ? ((8'hbe) == (8'hbf)) : (-(7'h48))), ((^(8'hac)) ? ((8'ha5) >= (8'ha3)) : (8'hba))} : (~^((~|(8'h9d)) ? ((8'ha2) ? (7'h40) : (8'had)) : ((7'h46) != (7'h46)))))))
(y, clk, wire425, wire424, wire423, wire422, wire421);
  output wire [(32'h7a0):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(2'h3):(1'h0)] wire425;
  input wire signed [(3'h5):(1'h0)] wire424;
  input wire [(4'hd):(1'h0)] wire423;
  input wire signed [(5'h10):(1'h0)] wire422;
  input wire signed [(5'h12):(1'h0)] wire421;
  wire [(4'hb):(1'h0)] wire570;
  wire [(5'h12):(1'h0)] wire532;
  wire [(5'h15):(1'h0)] wire530;
  wire signed [(3'h7):(1'h0)] wire529;
  wire [(5'h15):(1'h0)] wire528;
  wire signed [(4'h8):(1'h0)] wire512;
  wire signed [(5'h12):(1'h0)] wire511;
  wire [(4'hd):(1'h0)] wire510;
  wire [(5'h12):(1'h0)] wire506;
  wire [(5'h10):(1'h0)] wire480;
  wire signed [(4'h9):(1'h0)] wire427;
  wire signed [(4'ha):(1'h0)] wire426;
  reg signed [(4'h9):(1'h0)] reg573 = (1'h0);
  reg [(5'h12):(1'h0)] reg569 = (1'h0);
  reg [(4'hb):(1'h0)] reg567 = (1'h0);
  reg [(5'h11):(1'h0)] reg566 = (1'h0);
  reg [(5'h17):(1'h0)] reg562 = (1'h0);
  reg [(3'h7):(1'h0)] reg561 = (1'h0);
  reg [(5'h10):(1'h0)] reg558 = (1'h0);
  reg [(5'h12):(1'h0)] reg556 = (1'h0);
  reg [(5'h17):(1'h0)] reg554 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg552 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg551 = (1'h0);
  reg [(5'h11):(1'h0)] reg550 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg547 = (1'h0);
  reg [(5'h16):(1'h0)] reg546 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg542 = (1'h0);
  reg [(3'h6):(1'h0)] reg541 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg538 = (1'h0);
  reg [(4'hb):(1'h0)] reg537 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg534 = (1'h0);
  reg [(2'h2):(1'h0)] reg526 = (1'h0);
  reg [(3'h6):(1'h0)] reg524 = (1'h0);
  reg [(4'h9):(1'h0)] reg522 = (1'h0);
  reg [(3'h5):(1'h0)] reg520 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg519 = (1'h0);
  reg [(4'h9):(1'h0)] reg517 = (1'h0);
  reg [(3'h4):(1'h0)] reg515 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg513 = (1'h0);
  reg [(4'h9):(1'h0)] reg509 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg508 = (1'h0);
  reg [(5'h16):(1'h0)] reg507 = (1'h0);
  reg [(4'h9):(1'h0)] reg501 = (1'h0);
  reg [(4'ha):(1'h0)] reg498 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg495 = (1'h0);
  reg [(4'h8):(1'h0)] reg492 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg490 = (1'h0);
  reg [(4'hc):(1'h0)] reg489 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg486 = (1'h0);
  reg [(5'h10):(1'h0)] reg481 = (1'h0);
  reg [(5'h14):(1'h0)] reg476 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg474 = (1'h0);
  reg [(3'h7):(1'h0)] reg473 = (1'h0);
  reg [(4'hb):(1'h0)] reg470 = (1'h0);
  reg [(5'h10):(1'h0)] reg469 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg467 = (1'h0);
  reg [(5'h17):(1'h0)] reg453 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg463 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg460 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg454 = (1'h0);
  reg [(3'h4):(1'h0)] reg451 = (1'h0);
  reg [(4'hb):(1'h0)] reg449 = (1'h0);
  reg [(4'he):(1'h0)] reg446 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg445 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg444 = (1'h0);
  reg [(5'h14):(1'h0)] reg429 = (1'h0);
  reg [(4'hf):(1'h0)] reg443 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg442 = (1'h0);
  reg [(5'h11):(1'h0)] reg439 = (1'h0);
  reg [(3'h4):(1'h0)] reg435 = (1'h0);
  reg [(5'h18):(1'h0)] reg432 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg572 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg571 = (1'h0);
  reg [(4'h8):(1'h0)] reg568 = (1'h0);
  reg [(5'h11):(1'h0)] forvar565 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg564 = (1'h0);
  reg [(3'h5):(1'h0)] reg563 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg560 = (1'h0);
  reg signed [(4'he):(1'h0)] reg559 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg557 = (1'h0);
  reg [(2'h3):(1'h0)] reg555 = (1'h0);
  reg [(5'h15):(1'h0)] reg553 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar549 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg548 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg539 = (1'h0);
  reg [(4'ha):(1'h0)] reg545 = (1'h0);
  reg [(5'h16):(1'h0)] reg544 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg543 = (1'h0);
  reg [(2'h2):(1'h0)] reg540 = (1'h0);
  reg [(3'h5):(1'h0)] forvar539 = (1'h0);
  reg [(5'h14):(1'h0)] reg536 = (1'h0);
  reg [(5'h10):(1'h0)] reg535 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar533 = (1'h0);
  reg [(3'h4):(1'h0)] reg531 = (1'h0);
  reg [(4'ha):(1'h0)] reg527 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg525 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg523 = (1'h0);
  reg [(4'hf):(1'h0)] reg521 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg518 = (1'h0);
  reg [(4'hf):(1'h0)] reg516 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg514 = (1'h0);
  reg [(5'h10):(1'h0)] reg505 = (1'h0);
  reg [(4'he):(1'h0)] reg504 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg503 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg502 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg500 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg499 = (1'h0);
  reg [(4'h9):(1'h0)] forvar497 = (1'h0);
  reg [(3'h5):(1'h0)] reg496 = (1'h0);
  reg [(3'h6):(1'h0)] forvar494 = (1'h0);
  reg [(4'hf):(1'h0)] reg493 = (1'h0);
  reg [(2'h2):(1'h0)] reg491 = (1'h0);
  reg [(4'h9):(1'h0)] forvar488 = (1'h0);
  reg [(4'hb):(1'h0)] reg487 = (1'h0);
  reg [(4'hb):(1'h0)] reg485 = (1'h0);
  reg [(3'h4):(1'h0)] forvar484 = (1'h0);
  reg [(4'hc):(1'h0)] reg483 = (1'h0);
  reg [(3'h5):(1'h0)] forvar482 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg479 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar478 = (1'h0);
  reg [(3'h5):(1'h0)] reg477 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg475 = (1'h0);
  reg [(3'h5):(1'h0)] reg472 = (1'h0);
  reg [(4'hb):(1'h0)] reg471 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg468 = (1'h0);
  reg [(4'ha):(1'h0)] forvar466 = (1'h0);
  reg [(4'h9):(1'h0)] forvar447 = (1'h0);
  reg [(4'he):(1'h0)] forvar445 = (1'h0);
  reg [(5'h18):(1'h0)] reg465 = (1'h0);
  reg [(3'h6):(1'h0)] reg464 = (1'h0);
  reg [(3'h7):(1'h0)] reg462 = (1'h0);
  reg [(4'hc):(1'h0)] forvar461 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg459 = (1'h0);
  reg [(4'hf):(1'h0)] reg458 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg457 = (1'h0);
  reg [(4'hc):(1'h0)] reg456 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg455 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar453 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg452 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg450 = (1'h0);
  reg [(3'h7):(1'h0)] reg448 = (1'h0);
  reg [(4'hf):(1'h0)] reg447 = (1'h0);
  reg [(3'h6):(1'h0)] forvar441 = (1'h0);
  reg [(5'h15):(1'h0)] reg440 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg438 = (1'h0);
  reg [(3'h7):(1'h0)] reg437 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg436 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar434 = (1'h0);
  reg [(5'h13):(1'h0)] reg433 = (1'h0);
  reg [(4'hc):(1'h0)] reg431 = (1'h0);
  reg [(3'h7):(1'h0)] reg430 = (1'h0);
  reg [(5'h17):(1'h0)] forvar429 = (1'h0);
  reg [(5'h12):(1'h0)] reg428 = (1'h0);
  assign y = {wire570,
                 wire532,
                 wire530,
                 wire529,
                 wire528,
                 wire512,
                 wire511,
                 wire510,
                 wire506,
                 wire480,
                 wire427,
                 wire426,
                 reg573,
                 reg569,
                 reg567,
                 reg566,
                 reg562,
                 reg561,
                 reg558,
                 reg556,
                 reg554,
                 reg552,
                 reg551,
                 reg550,
                 reg547,
                 reg546,
                 reg542,
                 reg541,
                 reg538,
                 reg537,
                 reg534,
                 reg526,
                 reg524,
                 reg522,
                 reg520,
                 reg519,
                 reg517,
                 reg515,
                 reg513,
                 reg509,
                 reg508,
                 reg507,
                 reg501,
                 reg498,
                 reg495,
                 reg492,
                 reg490,
                 reg489,
                 reg486,
                 reg481,
                 reg476,
                 reg474,
                 reg473,
                 reg470,
                 reg469,
                 reg467,
                 reg453,
                 reg463,
                 reg460,
                 reg454,
                 reg451,
                 reg449,
                 reg446,
                 reg445,
                 reg444,
                 reg429,
                 reg443,
                 reg442,
                 reg439,
                 reg435,
                 reg432,
                 reg572,
                 reg571,
                 reg568,
                 forvar565,
                 reg564,
                 reg563,
                 reg560,
                 reg559,
                 reg557,
                 reg555,
                 reg553,
                 forvar549,
                 reg548,
                 reg539,
                 reg545,
                 reg544,
                 reg543,
                 reg540,
                 forvar539,
                 reg536,
                 reg535,
                 forvar533,
                 reg531,
                 reg527,
                 reg525,
                 reg523,
                 reg521,
                 reg518,
                 reg516,
                 reg514,
                 reg505,
                 reg504,
                 reg503,
                 reg502,
                 reg500,
                 reg499,
                 forvar497,
                 reg496,
                 forvar494,
                 reg493,
                 reg491,
                 forvar488,
                 reg487,
                 reg485,
                 forvar484,
                 reg483,
                 forvar482,
                 reg479,
                 forvar478,
                 reg477,
                 reg475,
                 reg472,
                 reg471,
                 reg468,
                 forvar466,
                 forvar447,
                 forvar445,
                 reg465,
                 reg464,
                 reg462,
                 forvar461,
                 reg459,
                 reg458,
                 reg457,
                 reg456,
                 reg455,
                 forvar453,
                 reg452,
                 reg450,
                 reg448,
                 reg447,
                 forvar441,
                 reg440,
                 reg438,
                 reg437,
                 reg436,
                 forvar434,
                 reg433,
                 reg431,
                 reg430,
                 forvar429,
                 reg428,
                 (1'h0)};
  assign wire426 = wire423[(1'h0):(1'h0)];
  assign wire427 = ($unsigned(((wire425 >>> (~&wire422)) ^ ((&wire424) - $unsigned(wire423)))) ?
                       wire425[(2'h2):(2'h2)] : wire426);
  always
    @(posedge clk) begin
      if ((^(wire426 == $unsigned((wire426[(3'h7):(3'h6)] ?
          {(8'h9d), wire427} : $unsigned(wire421))))))
        begin
          reg428 = wire423[(3'h6):(1'h0)];
          for (forvar429 = (1'h0); (forvar429 < (2'h3)); forvar429 = (forvar429 + (1'h1)))
            begin
              reg430 = $unsigned(wire427);
              reg431 = ($signed((wire421[(5'h10):(3'h6)] != $unsigned(wire423))) ?
                  ({(~wire427)} >= reg428) : (wire424[(1'h1):(1'h1)] <<< $signed(((~&wire424) ?
                      (wire423 ? (8'ha1) : (8'ha3)) : $unsigned(reg428)))));
              reg432 <= wire422[(3'h6):(1'h1)];
              reg433 = $unsigned((^~($signed(forvar429) ?
                  (wire427 < $signed(wire427)) : ((wire423 <= (8'hbb)) ?
                      forvar429 : (forvar429 ? reg432 : wire426)))));
            end
          for (forvar434 = (1'h0); (forvar434 < (1'h0)); forvar434 = (forvar434 + (1'h1)))
            begin
              reg435 <= ({$signed((wire424 * $unsigned(wire423)))} ?
                  wire427[(2'h3):(1'h0)] : $signed(reg428));
              reg436 = forvar434[(1'h1):(1'h1)];
              reg437 = (wire423 ?
                  (wire427 ~^ ($signed({forvar429, wire421}) ?
                      ((wire424 & forvar429) ?
                          reg430 : (reg436 < reg428)) : ((8'hba) ?
                          (wire422 ?
                              reg432 : (8'hb0)) : (~|reg435)))) : (^reg431[(3'h6):(3'h4)]));
              reg438 = (~$unsigned(reg431[(4'hb):(3'h7)]));
              reg439 <= $signed((wire425[(2'h2):(1'h1)] ?
                  (~((8'hbb) ^ wire421[(2'h3):(1'h0)])) : ($unsigned((|(8'hb7))) ?
                      (-(reg431 || wire423)) : (wire421 ?
                          $unsigned(forvar434) : $signed(forvar434)))));
            end
          reg440 = (reg428[(4'hf):(3'h4)] ?
              $unsigned((~($unsigned(wire427) ?
                  reg431 : reg438[(3'h7):(1'h1)]))) : ((&(|forvar429)) ?
                  forvar429[(4'hc):(1'h1)] : reg430));
          for (forvar441 = (1'h0); (forvar441 < (1'h1)); forvar441 = (forvar441 + (1'h1)))
            begin
              reg442 <= ($signed(((8'hba) ?
                      ($unsigned((8'hbc)) == $unsigned(reg436)) : wire426[(3'h6):(3'h5)])) ?
                  {reg433[(5'h12):(4'he)]} : wire421[(4'h9):(1'h0)]);
              reg443 <= forvar441[(3'h6):(1'h1)];
            end
        end
      else
        begin
          reg429 <= ((8'hb7) ?
              ((reg440[(4'h9):(1'h0)] ?
                  (forvar429[(3'h5):(3'h4)] >>> (reg442 ?
                      forvar434 : wire423)) : wire424) < (reg437[(3'h4):(1'h0)] ?
                  ((reg430 ? reg431 : reg428) ?
                      wire423[(3'h7):(2'h3)] : (reg443 < reg433)) : $unsigned((forvar434 ?
                      forvar434 : wire425)))) : wire422);
        end
      if (forvar429)
        begin
          if (($signed((^reg440)) ~^ reg435))
            begin
              reg444 <= (((|$signed($unsigned(wire424))) >>> (^reg442[(4'h9):(4'h9)])) ?
                  $unsigned({wire422, {forvar434}}) : {reg432,
                      forvar441[(3'h6):(2'h2)]});
              reg445 <= {{reg440,
                      $signed($signed((reg432 ? wire426 : (8'ha7))))}};
              reg446 <= forvar429[(4'ha):(3'h5)];
              reg447 = ($signed(wire425) ?
                  (~|(($signed((8'hbd)) || (reg436 ^~ reg432)) > {reg430,
                      (8'hb0)})) : {(|($signed(forvar441) ?
                          {reg435} : $signed(reg433))),
                      reg429});
              reg448 = $unsigned({$signed(((8'haa) ?
                      reg429[(4'hc):(2'h3)] : (reg439 || reg439)))});
            end
          else
            begin
              reg447 = {{$unsigned({(reg432 ? reg432 : (8'hb0)),
                          $unsigned(wire426)}),
                      {(!(+reg430))}},
                  ($signed((^~forvar441)) ?
                      (($signed(reg440) ? (reg446 ~^ reg443) : reg440) ?
                          ((8'had) && $unsigned((8'hb4))) : $unsigned(((8'ha7) ?
                              reg439 : (7'h45)))) : (^(~^(~(8'hb8)))))};
              reg449 <= (|(^(!$signed((-(7'h40))))));
              reg450 = $unsigned(((!$unsigned(reg428[(2'h2):(1'h1)])) <= reg432));
              reg451 <= ((reg433 >= $unsigned($unsigned(reg428))) ?
                  (!$unsigned(((reg450 ? reg428 : reg446) ?
                      (reg432 << reg449) : $signed(reg442)))) : {{reg432},
                      reg429[(4'hd):(4'h8)]});
              reg452 = ((&wire424) | $signed(((reg442 ?
                  forvar429[(4'hf):(4'hd)] : reg446) != ((reg428 ?
                  reg437 : reg437) * {reg439}))));
            end
          for (forvar453 = (1'h0); (forvar453 < (2'h3)); forvar453 = (forvar453 + (1'h1)))
            begin
              reg454 <= ($signed($signed($signed((reg445 + reg436)))) - reg450[(3'h5):(2'h2)]);
              reg455 = $unsigned($signed($signed($signed(reg437[(2'h3):(2'h3)]))));
              reg456 = reg454[(1'h0):(1'h0)];
            end
          reg457 = ({$unsigned(((wire423 ? reg430 : reg443) ?
                      reg439 : $signed(reg450))),
                  (forvar453[(4'h8):(1'h1)] ?
                      (reg431 ?
                          $unsigned(reg437) : $signed(forvar434)) : $unsigned($signed(reg429)))} ?
              (|reg432[(4'hc):(2'h2)]) : ((~{(^~reg444)}) ?
                  (-{reg437[(3'h6):(3'h5)]}) : $signed(((!reg439) ?
                      $signed((8'hb1)) : $unsigned((7'h45))))));
          if ($signed({(!{$unsigned(forvar453), (~&reg438)}),
              $unsigned((~^(!reg428)))}))
            begin
              reg458 = (reg446[(4'hb):(3'h5)] ?
                  $unsigned($signed($signed((wire421 < reg436)))) : (!((+$signed(reg456)) & $signed($signed(reg435)))));
              reg459 = {(-reg450)};
              reg460 <= (+reg435);
            end
          else
            begin
              reg458 = wire426[(3'h5):(3'h4)];
            end
          for (forvar461 = (1'h0); (forvar461 < (3'h4)); forvar461 = (forvar461 + (1'h1)))
            begin
              reg462 = (reg442[(4'h9):(4'h8)] ?
                  (^~((reg436 == (reg432 && reg444)) ?
                      (~^(reg457 ^ wire425)) : (&reg444))) : reg450);
              reg463 <= wire422[(4'h9):(1'h0)];
              reg464 = (reg437 ?
                  $signed(reg448[(3'h5):(2'h2)]) : $unsigned($signed(((forvar441 ?
                          reg442 : reg448) ?
                      (8'ha2) : (~|(8'hb8))))));
              reg465 = (reg443[(3'h6):(2'h3)] ?
                  $unsigned(({$signed(reg459), {reg443}} ?
                      (reg429 < reg429[(5'h11):(4'h9)]) : (^(~^reg428)))) : {forvar441[(3'h5):(2'h3)]});
            end
        end
      else
        begin
          if (((~reg448) ?
              ((8'hb0) ? reg429 : $signed(reg460[(5'h14):(1'h1)])) : (reg450 ?
                  ((^~(reg444 != reg446)) != $unsigned($signed(forvar461))) : ($signed(reg459) ?
                      reg463[(3'h6):(3'h4)] : reg465))))
            begin
              reg444 <= $unsigned(reg458[(4'ha):(4'h9)]);
            end
          else
            begin
              reg444 <= reg448[(2'h3):(2'h3)];
            end
          for (forvar445 = (1'h0); (forvar445 < (3'h4)); forvar445 = (forvar445 + (1'h1)))
            begin
              reg446 <= {((7'h40) ?
                      ((reg464[(1'h1):(1'h0)] ?
                              (reg462 + reg433) : $signed(wire424)) ?
                          reg436[(3'h4):(2'h3)] : $signed((~reg431))) : reg465[(3'h6):(1'h1)])};
            end
          for (forvar447 = (1'h0); (forvar447 < (1'h0)); forvar447 = (forvar447 + (1'h1)))
            begin
              reg449 <= (reg458 ?
                  ((^~(&$unsigned(reg456))) << (reg435 << (~(reg444 * reg451)))) : $unsigned((wire421 ?
                      $signed(forvar445) : $unsigned((~reg463)))));
              reg451 <= ($unsigned({reg458, (-$unsigned(reg456))}) ?
                  (~|((~&$signed(forvar441)) ?
                      (!$signed((8'hb6))) : $unsigned((forvar453 ?
                          reg443 : forvar453)))) : $unsigned(reg433[(1'h1):(1'h0)]));
              reg452 = {(reg465 ? (+wire425[(1'h0):(1'h0)]) : (|(8'hb6)))};
            end
          reg453 <= forvar445[(1'h1):(1'h0)];
          reg454 <= $unsigned((~&(~($unsigned(wire421) * reg450))));
        end
    end
  always
    @(posedge clk) begin
      for (forvar466 = (1'h0); (forvar466 < (2'h2)); forvar466 = (forvar466 + (1'h1)))
        begin
          reg467 <= ($signed($unsigned(reg451[(1'h0):(1'h0)])) ?
              reg446[(4'he):(4'hb)] : $signed((8'ha8)));
          if ((8'hb4))
            begin
              reg468 = reg449[(1'h1):(1'h0)];
            end
          else
            begin
              reg468 = ({((+wire422[(3'h5):(2'h2)]) < reg468),
                  reg432} >= ({{forvar466[(3'h7):(1'h1)],
                      ((8'hb1) ?
                          reg444 : wire427)}} || ($signed(reg439[(5'h11):(1'h0)]) ?
                  $unsigned(wire424) : (8'hac))));
              reg469 <= (-(~^(((~|forvar466) ?
                      (reg439 ^~ (8'ha0)) : (~wire427)) ?
                  forvar466[(4'ha):(4'ha)] : $unsigned($unsigned(reg445)))));
              reg470 <= ((|(reg460[(1'h1):(1'h1)] ?
                  reg449[(4'hb):(2'h3)] : $unsigned($unsigned((7'h4a))))) & $signed((reg460 ?
                  $signed(reg435) : reg469[(4'hd):(4'hb)])));
              reg471 = wire421[(2'h3):(1'h0)];
            end
          if (reg451[(1'h1):(1'h1)])
            begin
              reg472 = reg470;
              reg473 <= ((~|wire424[(1'h0):(1'h0)]) > wire424);
              reg474 <= $signed(($signed(reg432[(5'h14):(2'h3)]) ?
                  reg471 : forvar466[(1'h1):(1'h1)]));
              reg475 = reg432;
            end
          else
            begin
              reg472 = $signed(reg454);
              reg475 = $signed({reg454[(3'h6):(1'h1)]});
              reg476 <= ($unsigned((((reg453 ?
                          reg454 : reg470) >>> (reg475 * reg444)) ?
                      {{wire421},
                          (reg460 && wire422)} : ($signed(wire423) >> reg439[(2'h2):(2'h2)]))) ?
                  wire422[(1'h0):(1'h0)] : (~(reg473 < $signed($unsigned(reg432)))));
              reg477 = $signed({{$signed($unsigned(reg468))},
                  $signed(wire425)});
            end
          for (forvar478 = (1'h0); (forvar478 < (1'h0)); forvar478 = (forvar478 + (1'h1)))
            begin
              reg479 = (reg445 ? reg474 : $unsigned(reg449));
            end
        end
    end
  assign wire480 = $unsigned((^reg445[(3'h6):(1'h1)]));
  always
    @(posedge clk) begin
      reg481 <= reg442;
      for (forvar482 = (1'h0); (forvar482 < (2'h3)); forvar482 = (forvar482 + (1'h1)))
        begin
          reg483 = $signed(({((~^reg481) ?
                      (reg467 >= wire427) : (reg442 ? reg435 : wire480)),
                  $unsigned($signed((8'hbe)))} ?
              $signed($unsigned(reg435[(2'h2):(2'h2)])) : (wire425 ?
                  $signed(((7'h48) ?
                      reg432 : reg470)) : (^~$unsigned((8'ha4))))));
          for (forvar484 = (1'h0); (forvar484 < (1'h0)); forvar484 = (forvar484 + (1'h1)))
            begin
              reg485 = wire480[(4'hf):(4'h8)];
            end
          reg486 <= (8'hb0);
          reg487 = {reg467,
              ($signed((((8'hb2) + reg435) ?
                  (reg442 >= forvar482) : (reg432 == reg469))) > $signed($unsigned((reg443 >> reg470))))};
        end
      for (forvar488 = (1'h0); (forvar488 < (2'h3)); forvar488 = (forvar488 + (1'h1)))
        begin
          if (reg451[(1'h1):(1'h0)])
            begin
              reg489 <= reg451[(1'h1):(1'h1)];
              reg490 <= (((8'hb6) | (~(!(reg486 ?
                  (7'h43) : reg444)))) - ((8'hae) ~^ reg443));
            end
          else
            begin
              reg491 = (((~&(!$unsigned(reg470))) ^~ $unsigned($unsigned($unsigned(reg432)))) | $signed(reg435));
              reg492 <= $unsigned((reg449 ? reg445 : (&forvar482)));
              reg493 = $unsigned($unsigned($unsigned(reg476[(3'h7):(3'h7)])));
            end
          for (forvar494 = (1'h0); (forvar494 < (3'h4)); forvar494 = (forvar494 + (1'h1)))
            begin
              reg495 <= (|$signed((8'haf)));
              reg496 = (~&reg453);
            end
          for (forvar497 = (1'h0); (forvar497 < (2'h2)); forvar497 = (forvar497 + (1'h1)))
            begin
              reg498 <= reg442[(4'ha):(4'h8)];
              reg499 = $signed(forvar494);
              reg500 = $signed((^$unsigned(forvar484)));
              reg501 <= reg487;
              reg502 = $signed(reg473);
            end
          if (reg432)
            begin
              reg503 = (8'ha4);
              reg504 = (~((~forvar497[(1'h1):(1'h1)]) >> (reg503 ?
                  wire424 : reg469[(4'h9):(3'h6)])));
              reg505 = reg445[(4'he):(4'hd)];
            end
          else
            begin
              reg503 = $signed(reg496);
            end
        end
    end
  assign wire506 = ({{(~wire426[(4'h8):(1'h1)]), $unsigned({wire427})},
                           reg444[(4'he):(3'h5)]} ?
                       wire421 : reg474);
  always
    @(posedge clk) begin
      reg507 <= (reg443 ? (~reg489) : reg449);
      reg508 <= ($signed(($unsigned((reg467 == reg432)) < ((~reg444) - (^reg446)))) ?
          reg451[(1'h1):(1'h0)] : (($signed(reg446[(1'h0):(1'h0)]) == ((8'hb7) ?
              (^~reg446) : $signed(reg454))) == wire423));
    end
  always
    @(posedge clk) begin
      reg509 <= {reg498};
    end
  assign wire510 = reg467[(5'h18):(5'h15)];
  assign wire511 = wire480;
  assign wire512 = reg449;
  always
    @(posedge clk) begin
      if ({reg486[(4'he):(2'h2)]})
        begin
          reg513 <= (!$signed({(~&((7'h4a) ? reg449 : (7'h4a))),
              $unsigned($unsigned(reg439))}));
        end
      else
        begin
          reg514 = (-((^~((8'hae) & reg435)) ?
              (((^wire506) * (reg495 ?
                  reg435 : reg435)) == $signed((reg474 - reg490))) : wire480));
          reg515 <= ((~(~wire510)) - ((reg513[(3'h7):(2'h3)] * $unsigned(((8'h9c) ^ reg481))) ?
              reg467[(5'h17):(4'hf)] : wire480));
          if (((!(reg486[(3'h5):(3'h4)] ?
              (reg513[(3'h4):(1'h1)] ^~ (+wire421)) : ((^~wire512) ?
                  (reg507 <= reg429) : (wire426 ?
                      (8'h9f) : reg446)))) ^~ $signed(reg489[(3'h4):(3'h4)])))
            begin
              reg516 = (-$signed($signed($unsigned($signed(reg509)))));
              reg517 <= $signed($unsigned(($signed(reg445[(5'h14):(5'h11)]) ?
                  $unsigned(reg470) : (wire506 >= (^~reg515)))));
              reg518 = (|reg501);
              reg519 <= ((^$unsigned(reg449[(2'h2):(1'h0)])) >>> ($signed($signed(reg429)) ?
                  $signed({reg443[(4'ha):(1'h0)]}) : reg492[(1'h0):(1'h0)]));
              reg520 <= {{reg444}};
            end
          else
            begin
              reg517 <= reg492;
              reg518 = $unsigned((reg520 ~^ ({(wire426 ? (8'hb4) : reg513)} ?
                  reg443[(4'h8):(1'h0)] : ($signed((8'hb2)) ?
                      (reg444 ? reg445 : wire480) : {reg449}))));
              reg521 = ({reg501,
                      ($signed({reg490}) ?
                          $signed((~|reg443)) : ((8'h9f) ?
                              (wire422 * wire511) : (!reg432)))} ?
                  reg515 : reg467[(5'h12):(5'h12)]);
              reg522 <= (~^reg463[(4'h8):(3'h5)]);
            end
          reg523 = reg444;
          reg524 <= reg439;
        end
      if ($unsigned($unsigned((((reg490 >= reg473) != (~|(8'ha9))) ?
          ((~wire506) ?
              ((8'hb2) ?
                  wire425 : reg446) : (-reg467)) : $unsigned(wire423[(4'h8):(1'h1)])))))
        begin
          reg525 = reg509[(4'h9):(1'h1)];
          reg526 <= $unsigned((reg460[(4'h8):(3'h5)] - $signed((~^(reg470 ?
              (8'hb7) : (8'hb6))))));
          reg527 = ($unsigned((7'h42)) ? reg516 : (8'hb0));
        end
      else
        begin
          reg525 = (8'ha1);
        end
    end
  assign wire528 = ($signed(((~&{reg463, reg463}) ?
                       $signed($signed(reg449)) : reg517[(4'h9):(4'h8)])) >> ($unsigned($unsigned(((8'hb2) ?
                           reg473 : reg439))) ?
                       $unsigned(((reg467 | reg526) != reg451[(2'h3):(1'h1)])) : $signed($unsigned($signed(wire423)))));
  assign wire529 = $signed({{(8'hbc)},
                       (wire528 ? (-(-reg470)) : $unsigned(reg449))});
  assign wire530 = (($signed((((8'hb9) ? wire424 : wire424) ?
                       (8'ha1) : $unsigned(reg517))) == {reg473[(2'h2):(1'h0)]}) == wire427[(3'h7):(2'h3)]);
  always
    @(posedge clk) begin
      reg531 = $unsigned(((^~$signed({reg515, reg445})) ?
          {((reg486 || reg449) ?
                  ((8'hbe) ?
                      reg453 : reg524) : (reg486 && reg435))} : {(~wire427)}));
    end
  assign wire532 = {reg517[(3'h4):(3'h4)], reg486};
  always
    @(posedge clk) begin
      for (forvar533 = (1'h0); (forvar533 < (1'h0)); forvar533 = (forvar533 + (1'h1)))
        begin
          reg534 <= reg513;
          reg535 = reg463;
        end
    end
  always
    @(posedge clk) begin
      reg536 = ((((reg489[(1'h1):(1'h0)] ? (wire512 <= reg446) : reg473) ?
                  {((7'h41) ? wire425 : wire480)} : reg520) ?
              reg501[(1'h0):(1'h0)] : $signed($signed($signed(wire506)))) ?
          ($unsigned({$signed(reg453)}) >> ((7'h43) & (8'ha5))) : reg490[(3'h7):(1'h0)]);
      if ((8'haf))
        begin
          reg537 <= $unsigned((~(((&reg517) ~^ (+reg520)) & (reg460[(5'h16):(4'ha)] >= (~^reg460)))));
          reg538 <= {(~^reg492[(1'h0):(1'h0)]),
              $unsigned(wire511[(4'hc):(4'hb)])};
          for (forvar539 = (1'h0); (forvar539 < (2'h3)); forvar539 = (forvar539 + (1'h1)))
            begin
              reg540 = $signed(wire423[(4'hd):(2'h2)]);
              reg541 <= (-reg460);
              reg542 <= ($unsigned(reg522[(1'h0):(1'h0)]) ?
                  ((7'h42) + ((reg453 ?
                      (wire422 ? reg481 : reg486) : (~^reg476)) ^~ {(reg444 ?
                          wire423 : reg486),
                      (wire480 >>> wire421)})) : (wire421 ?
                      {(^reg444[(3'h6):(3'h5)]), (7'h44)} : wire532));
            end
          if ($unsigned($unsigned(($signed($signed(reg508)) ?
              ((wire425 ? reg445 : (7'h49)) != (reg486 ?
                  wire528 : reg429)) : reg538))))
            begin
              reg543 = (reg524[(2'h3):(2'h3)] < reg524);
              reg544 = ($signed($unsigned($signed(reg522))) >= $unsigned(((reg446[(2'h2):(1'h0)] ?
                      $unsigned(reg536) : {reg541}) ?
                  (reg474 <= (8'haa)) : ({forvar539} ~^ {reg534, reg476}))));
              reg545 = ((^~({$unsigned(reg536), (reg432 ^ (8'hae))} ?
                      ((reg543 && reg442) ?
                          wire506[(4'hb):(4'h9)] : (reg541 > forvar539)) : ($unsigned(reg524) >= wire529[(2'h3):(1'h0)]))) ?
                  {reg517} : (!((&reg451) & ({wire506,
                      wire427} | (~^reg476)))));
            end
          else
            begin
              reg546 <= ($signed($unsigned($unsigned((reg463 < reg432)))) ?
                  ($unsigned($unsigned(((7'h42) ? reg469 : (7'h40)))) ?
                      $unsigned(reg444) : (^$unsigned($signed((8'h9d))))) : $unsigned((((reg470 ?
                      reg492 : reg537) >> $signed(reg542)) > $signed((reg463 ?
                      (8'ha3) : (8'ha1))))));
              reg547 <= reg538;
            end
        end
      else
        begin
          if ((&$signed(({$signed(reg474), $unsigned(reg454)} ?
              {{wire422}} : ($unsigned((8'ha8)) ?
                  reg542 : $unsigned(reg544))))))
            begin
              reg539 = reg474;
              reg541 <= $unsigned(reg513);
              reg542 <= ($unsigned(wire530) | wire427);
              reg546 <= (~|({$signed((wire422 ? reg539 : reg432))} ?
                  {$signed((^~reg429))} : $signed($unsigned($signed(wire421)))));
              reg548 = {((reg432 ?
                      $unsigned(reg470[(3'h4):(1'h0)]) : reg470[(4'hb):(2'h3)]) - ($unsigned($unsigned(wire480)) <= $unsigned(reg544[(4'hc):(2'h3)])))};
            end
          else
            begin
              reg537 <= wire529;
            end
          for (forvar549 = (1'h0); (forvar549 < (2'h2)); forvar549 = (forvar549 + (1'h1)))
            begin
              reg550 <= $signed((((~|(^~reg444)) >> $unsigned($signed(reg508))) ?
                  $unsigned(((reg490 ? reg544 : reg522) ?
                      $signed(forvar539) : (~&wire423))) : (&reg507[(2'h3):(1'h0)])));
              reg551 <= (~|wire511);
            end
          if (reg545)
            begin
              reg552 <= $unsigned($unsigned($signed(((reg537 ?
                      reg492 : (8'hac)) ?
                  $unsigned(reg542) : $signed(reg541)))));
            end
          else
            begin
              reg553 = $signed((($signed($unsigned(wire506)) ^~ $signed((7'h47))) && wire422[(2'h2):(1'h0)]));
              reg554 <= $signed({(reg547 <<< $unsigned({forvar549, reg519}))});
              reg555 = {($unsigned(reg474[(4'hc):(2'h2)]) ?
                      ((reg546 ~^ (wire511 ? reg481 : reg536)) ?
                          (+(+wire529)) : (~|(reg446 ?
                              reg554 : reg498))) : ((reg507[(5'h14):(4'hc)] | (reg513 ?
                              reg432 : reg540)) ?
                          $signed((~(8'ha3))) : (8'ha9))),
                  reg463[(4'ha):(4'h9)]};
              reg556 <= ($signed((~^reg449[(4'h9):(4'h8)])) >= ($signed($signed(((8'hb2) ?
                      wire425 : reg513))) ?
                  (wire530[(3'h5):(3'h4)] ?
                      (~|wire530) : reg467[(2'h3):(1'h0)]) : $unsigned($unsigned(reg501))));
            end
        end
      reg557 = ((8'h9f) >> reg446);
      if ($unsigned($unsigned($signed(wire530))))
        begin
          if ((($unsigned(({reg517, (8'hb6)} ?
              $unsigned(reg548) : reg545[(3'h6):(1'h1)])) ~^ $unsigned($signed($unsigned(reg435)))) < {($signed((-reg547)) > $signed(reg515)),
              reg446[(4'hd):(4'hd)]}))
            begin
              reg558 <= $signed((|reg542[(1'h0):(1'h0)]));
              reg559 = reg539[(4'h8):(1'h0)];
            end
          else
            begin
              reg558 <= $signed(reg446[(3'h4):(2'h3)]);
              reg559 = reg489;
            end
        end
      else
        begin
          if ($signed(((&{$unsigned(reg517)}) ?
              (|(8'ha3)) : reg556[(3'h5):(2'h3)])))
            begin
              reg558 <= wire529[(2'h3):(2'h2)];
            end
          else
            begin
              reg559 = ((reg507[(5'h15):(5'h11)] > reg498[(1'h1):(1'h0)]) - {reg547[(5'h14):(1'h1)]});
              reg560 = wire511[(3'h7):(3'h5)];
              reg561 <= reg557;
              reg562 <= $signed(wire422[(4'h9):(3'h6)]);
              reg563 = {reg538};
            end
          reg564 = (~^reg555);
          for (forvar565 = (1'h0); (forvar565 < (1'h1)); forvar565 = (forvar565 + (1'h1)))
            begin
              reg566 <= forvar549;
              reg567 <= $unsigned((((reg537[(4'ha):(4'ha)] <<< $signed(reg515)) ?
                  $signed({reg509, reg524}) : reg526) ^ reg566[(4'hd):(3'h6)]));
            end
          reg568 = {reg550};
          if ({(-(reg547 <<< reg546))})
            begin
              reg569 <= (!($signed($signed($unsigned((8'ha6)))) >>> $signed(((wire424 - reg470) == ((8'hb8) ?
                  reg492 : (8'hb1))))));
            end
          else
            begin
              reg569 <= $unsigned(($unsigned(wire506[(5'h10):(4'h9)]) ?
                  (~($unsigned(reg520) || (~^reg517))) : wire512));
            end
        end
    end
  assign wire570 = (-reg495);
  always
    @(posedge clk) begin
      reg571 = (&(({reg515,
          (~^wire424)} << reg517[(2'h2):(2'h2)]) && ($unsigned($unsigned(reg498)) != $unsigned((8'hb6)))));
      reg572 = ((reg534[(1'h1):(1'h0)] ?
          reg569[(5'h12):(4'ha)] : reg558[(2'h2):(1'h1)]) == $unsigned(($unsigned((wire570 ?
              reg561 : wire532)) ?
          $unsigned((wire422 ? reg524 : (8'hbd))) : reg508[(1'h0):(1'h0)])));
      reg573 <= ($signed(wire424[(2'h3):(1'h1)]) ?
          reg547 : (~|{wire512[(3'h6):(2'h3)], (|reg460)}));
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module962
#(parameter param1163 = ((8'ha2) >= ((((+(8'hac)) & ((7'h49) ? (8'h9d) : (7'h42))) ? (((8'hab) ? (8'hbd) : (7'h47)) <= {(7'h40), (8'ha8)}) : (8'hb6)) ? (8'hbb) : (({(8'ha9), (8'ha8)} ^ (~^(8'hbb))) ? (-((7'h47) ^ (8'ha7))) : (7'h48)))))
(y, clk, wire966, wire965, wire964, wire963);
  output wire [(32'had3):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire [(4'hd):(1'h0)] wire966;
  input wire [(2'h2):(1'h0)] wire965;
  input wire [(4'hc):(1'h0)] wire964;
  input wire signed [(4'hd):(1'h0)] wire963;
  wire [(5'h12):(1'h0)] wire1142;
  wire signed [(5'h12):(1'h0)] wire1141;
  wire signed [(4'hc):(1'h0)] wire1140;
  wire [(4'ha):(1'h0)] wire1139;
  wire signed [(5'h11):(1'h0)] wire1122;
  wire signed [(5'h14):(1'h0)] wire1103;
  wire [(4'h8):(1'h0)] wire1056;
  wire signed [(4'h9):(1'h0)] wire996;
  wire [(5'h10):(1'h0)] wire995;
  wire [(3'h5):(1'h0)] wire994;
  wire [(5'h15):(1'h0)] wire993;
  reg signed [(2'h3):(1'h0)] reg1162 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1161 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1159 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg1158 = (1'h0);
  reg [(4'ha):(1'h0)] reg1157 = (1'h0);
  reg [(5'h17):(1'h0)] reg1155 = (1'h0);
  reg [(3'h7):(1'h0)] reg1153 = (1'h0);
  reg [(4'ha):(1'h0)] reg1152 = (1'h0);
  reg [(4'h8):(1'h0)] reg1149 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1147 = (1'h0);
  reg [(4'hd):(1'h0)] reg1138 = (1'h0);
  reg [(5'h13):(1'h0)] reg1132 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1127 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1126 = (1'h0);
  reg [(4'h9):(1'h0)] reg1125 = (1'h0);
  reg [(3'h4):(1'h0)] reg1124 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1120 = (1'h0);
  reg [(2'h2):(1'h0)] reg1119 = (1'h0);
  reg [(2'h2):(1'h0)] reg1118 = (1'h0);
  reg [(5'h15):(1'h0)] reg1117 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1116 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1113 = (1'h0);
  reg [(3'h7):(1'h0)] reg1112 = (1'h0);
  reg [(5'h13):(1'h0)] reg1111 = (1'h0);
  reg [(2'h3):(1'h0)] reg1109 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1108 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1105 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1099 = (1'h0);
  reg [(3'h7):(1'h0)] reg1093 = (1'h0);
  reg [(3'h7):(1'h0)] reg1091 = (1'h0);
  reg [(2'h3):(1'h0)] reg1090 = (1'h0);
  reg [(4'he):(1'h0)] reg1088 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1087 = (1'h0);
  reg [(5'h15):(1'h0)] reg1085 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1084 = (1'h0);
  reg [(5'h17):(1'h0)] reg1082 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1080 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1078 = (1'h0);
  reg [(2'h3):(1'h0)] reg1075 = (1'h0);
  reg [(5'h12):(1'h0)] reg1074 = (1'h0);
  reg [(5'h12):(1'h0)] reg1073 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1072 = (1'h0);
  reg [(4'h9):(1'h0)] reg1070 = (1'h0);
  reg [(3'h5):(1'h0)] reg1067 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1055 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg1053 = (1'h0);
  reg [(5'h12):(1'h0)] reg1050 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1048 = (1'h0);
  reg [(3'h6):(1'h0)] reg1040 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg1045 = (1'h0);
  reg [(5'h11):(1'h0)] reg1043 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg1042 = (1'h0);
  reg signed [(4'he):(1'h0)] reg1038 = (1'h0);
  reg [(5'h12):(1'h0)] reg1037 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg1036 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1035 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1033 = (1'h0);
  reg [(5'h11):(1'h0)] reg1030 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1028 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1026 = (1'h0);
  reg [(5'h11):(1'h0)] reg1024 = (1'h0);
  reg [(3'h4):(1'h0)] reg1021 = (1'h0);
  reg [(5'h17):(1'h0)] reg1020 = (1'h0);
  reg [(4'h8):(1'h0)] reg1016 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1015 = (1'h0);
  reg [(2'h3):(1'h0)] reg1013 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1012 = (1'h0);
  reg [(4'h8):(1'h0)] reg1002 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg998 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1010 = (1'h0);
  reg [(4'hd):(1'h0)] reg1009 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg1007 = (1'h0);
  reg [(4'hf):(1'h0)] reg1005 = (1'h0);
  reg [(4'h8):(1'h0)] reg1004 = (1'h0);
  reg [(4'h9):(1'h0)] reg999 = (1'h0);
  reg [(4'he):(1'h0)] reg997 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg992 = (1'h0);
  reg [(5'h13):(1'h0)] reg989 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg985 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg981 = (1'h0);
  reg [(4'hb):(1'h0)] reg979 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg977 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg975 = (1'h0);
  reg [(4'hd):(1'h0)] reg974 = (1'h0);
  reg [(3'h7):(1'h0)] reg973 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg972 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg970 = (1'h0);
  reg [(3'h5):(1'h0)] reg1160 = (1'h0);
  reg [(3'h6):(1'h0)] forvar1157 = (1'h0);
  reg [(5'h18):(1'h0)] reg1156 = (1'h0);
  reg [(5'h14):(1'h0)] reg1150 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1149 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1146 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1156 = (1'h0);
  reg [(4'h8):(1'h0)] reg1154 = (1'h0);
  reg [(5'h13):(1'h0)] reg1151 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1150 = (1'h0);
  reg [(4'h8):(1'h0)] reg1148 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar1146 = (1'h0);
  reg [(5'h14):(1'h0)] reg1145 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1144 = (1'h0);
  reg [(4'hd):(1'h0)] forvar1143 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1137 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1136 = (1'h0);
  reg [(3'h6):(1'h0)] reg1135 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1134 = (1'h0);
  reg [(2'h3):(1'h0)] reg1133 = (1'h0);
  reg [(4'hf):(1'h0)] forvar1131 = (1'h0);
  reg [(5'h13):(1'h0)] reg1130 = (1'h0);
  reg [(5'h15):(1'h0)] reg1129 = (1'h0);
  reg [(5'h17):(1'h0)] reg1128 = (1'h0);
  reg [(4'hc):(1'h0)] reg1123 = (1'h0);
  reg [(4'hc):(1'h0)] reg1121 = (1'h0);
  reg signed [(4'hc):(1'h0)] forvar1115 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1114 = (1'h0);
  reg [(5'h14):(1'h0)] reg1110 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1106 = (1'h0);
  reg [(4'he):(1'h0)] forvar1105 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg1107 = (1'h0);
  reg [(2'h3):(1'h0)] forvar1106 = (1'h0);
  reg [(4'hd):(1'h0)] reg1104 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg1102 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1101 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1100 = (1'h0);
  reg [(4'hb):(1'h0)] reg1098 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1097 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg1096 = (1'h0);
  reg [(4'he):(1'h0)] reg1095 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1094 = (1'h0);
  reg [(5'h10):(1'h0)] forvar1092 = (1'h0);
  reg [(5'h14):(1'h0)] reg1089 = (1'h0);
  reg [(3'h5):(1'h0)] reg1086 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar1083 = (1'h0);
  reg [(4'he):(1'h0)] reg1081 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg1079 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1077 = (1'h0);
  reg [(4'ha):(1'h0)] reg1071 = (1'h0);
  reg [(4'he):(1'h0)] reg1076 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1071 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg1069 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1068 = (1'h0);
  reg [(5'h15):(1'h0)] reg1057 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1066 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1065 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1064 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1063 = (1'h0);
  reg [(3'h4):(1'h0)] reg1062 = (1'h0);
  reg [(5'h14):(1'h0)] reg1061 = (1'h0);
  reg [(5'h12):(1'h0)] reg1060 = (1'h0);
  reg [(2'h2):(1'h0)] reg1059 = (1'h0);
  reg [(4'he):(1'h0)] reg1058 = (1'h0);
  reg [(4'hc):(1'h0)] forvar1057 = (1'h0);
  reg [(5'h11):(1'h0)] forvar1054 = (1'h0);
  reg [(5'h17):(1'h0)] reg1052 = (1'h0);
  reg [(4'he):(1'h0)] reg1051 = (1'h0);
  reg [(5'h13):(1'h0)] reg1049 = (1'h0);
  reg [(2'h2):(1'h0)] forvar1048 = (1'h0);
  reg [(5'h12):(1'h0)] reg1047 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1046 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar1041 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1044 = (1'h0);
  reg [(5'h15):(1'h0)] reg1041 = (1'h0);
  reg [(5'h15):(1'h0)] forvar1040 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg1039 = (1'h0);
  reg [(5'h10):(1'h0)] reg1034 = (1'h0);
  reg [(4'he):(1'h0)] reg1032 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg1031 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg1029 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg1027 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg1025 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg1023 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg1022 = (1'h0);
  reg [(5'h18):(1'h0)] reg1019 = (1'h0);
  reg [(5'h15):(1'h0)] reg1018 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg1017 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg1014 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar1011 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar997 = (1'h0);
  reg [(2'h2):(1'h0)] reg1008 = (1'h0);
  reg [(4'hf):(1'h0)] reg1006 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg1003 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar1002 = (1'h0);
  reg [(4'he):(1'h0)] reg1001 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg1000 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar998 = (1'h0);
  reg [(2'h3):(1'h0)] reg991 = (1'h0);
  reg [(4'hc):(1'h0)] reg990 = (1'h0);
  reg [(5'h10):(1'h0)] reg988 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg987 = (1'h0);
  reg [(3'h4):(1'h0)] reg986 = (1'h0);
  reg [(5'h15):(1'h0)] reg984 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar983 = (1'h0);
  reg [(5'h11):(1'h0)] reg982 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg980 = (1'h0);
  reg [(5'h18):(1'h0)] reg976 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg969 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg978 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar976 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg971 = (1'h0);
  reg [(4'ha):(1'h0)] forvar969 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg968 = (1'h0);
  reg [(3'h5):(1'h0)] reg967 = (1'h0);
  assign y = {wire1142,
                 wire1141,
                 wire1140,
                 wire1139,
                 wire1122,
                 wire1103,
                 wire1056,
                 wire996,
                 wire995,
                 wire994,
                 wire993,
                 reg1162,
                 reg1161,
                 reg1159,
                 reg1158,
                 reg1157,
                 reg1155,
                 reg1153,
                 reg1152,
                 reg1149,
                 reg1147,
                 reg1138,
                 reg1132,
                 reg1127,
                 reg1126,
                 reg1125,
                 reg1124,
                 reg1120,
                 reg1119,
                 reg1118,
                 reg1117,
                 reg1116,
                 reg1113,
                 reg1112,
                 reg1111,
                 reg1109,
                 reg1108,
                 reg1105,
                 reg1099,
                 reg1093,
                 reg1091,
                 reg1090,
                 reg1088,
                 reg1087,
                 reg1085,
                 reg1084,
                 reg1082,
                 reg1080,
                 reg1078,
                 reg1075,
                 reg1074,
                 reg1073,
                 reg1072,
                 reg1070,
                 reg1067,
                 reg1055,
                 reg1053,
                 reg1050,
                 reg1048,
                 reg1040,
                 reg1045,
                 reg1043,
                 reg1042,
                 reg1038,
                 reg1037,
                 reg1036,
                 reg1035,
                 reg1033,
                 reg1030,
                 reg1028,
                 reg1026,
                 reg1024,
                 reg1021,
                 reg1020,
                 reg1016,
                 reg1015,
                 reg1013,
                 reg1012,
                 reg1002,
                 reg998,
                 reg1010,
                 reg1009,
                 reg1007,
                 reg1005,
                 reg1004,
                 reg999,
                 reg997,
                 reg992,
                 reg989,
                 reg985,
                 reg981,
                 reg979,
                 reg977,
                 reg975,
                 reg974,
                 reg973,
                 reg972,
                 reg970,
                 reg1160,
                 forvar1157,
                 reg1156,
                 reg1150,
                 forvar1149,
                 reg1146,
                 forvar1156,
                 reg1154,
                 reg1151,
                 forvar1150,
                 reg1148,
                 forvar1146,
                 reg1145,
                 reg1144,
                 forvar1143,
                 reg1137,
                 reg1136,
                 reg1135,
                 reg1134,
                 reg1133,
                 forvar1131,
                 reg1130,
                 reg1129,
                 reg1128,
                 reg1123,
                 reg1121,
                 forvar1115,
                 reg1114,
                 reg1110,
                 reg1106,
                 forvar1105,
                 reg1107,
                 forvar1106,
                 reg1104,
                 reg1102,
                 reg1101,
                 reg1100,
                 reg1098,
                 reg1097,
                 reg1096,
                 reg1095,
                 reg1094,
                 forvar1092,
                 reg1089,
                 reg1086,
                 forvar1083,
                 reg1081,
                 reg1079,
                 reg1077,
                 reg1071,
                 reg1076,
                 forvar1071,
                 reg1069,
                 reg1068,
                 reg1057,
                 forvar1066,
                 reg1065,
                 reg1064,
                 reg1063,
                 reg1062,
                 reg1061,
                 reg1060,
                 reg1059,
                 reg1058,
                 forvar1057,
                 forvar1054,
                 reg1052,
                 reg1051,
                 reg1049,
                 forvar1048,
                 reg1047,
                 reg1046,
                 forvar1041,
                 reg1044,
                 reg1041,
                 forvar1040,
                 reg1039,
                 reg1034,
                 reg1032,
                 reg1031,
                 reg1029,
                 reg1027,
                 reg1025,
                 reg1023,
                 reg1022,
                 reg1019,
                 reg1018,
                 reg1017,
                 reg1014,
                 forvar1011,
                 forvar997,
                 reg1008,
                 reg1006,
                 reg1003,
                 forvar1002,
                 reg1001,
                 reg1000,
                 forvar998,
                 reg991,
                 reg990,
                 reg988,
                 reg987,
                 reg986,
                 reg984,
                 forvar983,
                 reg982,
                 reg980,
                 reg976,
                 reg969,
                 reg978,
                 forvar976,
                 reg971,
                 forvar969,
                 reg968,
                 reg967,
                 (1'h0)};
  always
    @(posedge clk) begin
      reg967 = (8'ha8);
      reg968 = wire965[(1'h0):(1'h0)];
      if (($unsigned(wire964[(4'ha):(4'ha)]) ? wire965 : (+wire966)))
        begin
          for (forvar969 = (1'h0); (forvar969 < (1'h0)); forvar969 = (forvar969 + (1'h1)))
            begin
              reg970 <= $signed($unsigned((~^((wire964 <<< wire965) ?
                  (~|reg967) : (reg968 ? reg968 : (8'ha8))))));
              reg971 = ((~(reg970 <<< forvar969)) == $signed(wire964[(4'h9):(1'h0)]));
            end
          if (forvar969)
            begin
              reg972 <= ((reg968[(4'hb):(3'h5)] ?
                      (((|forvar969) ?
                          (forvar969 ?
                              (8'ha0) : (7'h45)) : $signed((8'ha8))) && $signed($signed(reg970))) : {($signed(reg967) >= forvar969[(2'h2):(2'h2)])}) ?
                  (8'ha4) : wire965);
              reg973 <= $signed((8'hac));
              reg974 <= wire963;
            end
          else
            begin
              reg972 <= {$signed((~^$signed({(8'h9d), wire963})))};
              reg973 <= (&(~^wire965));
              reg974 <= forvar969[(3'h6):(1'h1)];
              reg975 <= ({(($unsigned(reg973) ?
                          (reg973 ?
                              wire965 : wire965) : $unsigned(reg967)) && $signed($signed(reg970))),
                      (wire964[(4'hb):(1'h1)] ?
                          (^{(8'ha7)}) : ($signed(reg968) >= (reg968 ?
                              reg973 : reg967)))} ?
                  (8'hb3) : $unsigned(reg974));
            end
          for (forvar976 = (1'h0); (forvar976 < (1'h0)); forvar976 = (forvar976 + (1'h1)))
            begin
              reg977 <= (|(reg968[(1'h0):(1'h0)] <<< (~|$signed((reg975 ^ wire963)))));
              reg978 = (reg972 ? (8'hb0) : (8'h9d));
            end
          reg979 <= $signed(wire966[(3'h4):(3'h4)]);
        end
      else
        begin
          if (((($unsigned({reg970}) * forvar969[(1'h0):(1'h0)]) || forvar976[(2'h2):(2'h2)]) ?
              (|(reg974 ?
                  $signed((|wire966)) : (~^((8'ha0) >>> reg968)))) : (&(~^$signed(reg970[(4'hf):(3'h4)])))))
            begin
              reg969 = $signed({$unsigned(forvar976[(1'h1):(1'h0)]), reg972});
            end
          else
            begin
              reg969 = reg977[(2'h2):(1'h1)];
              reg971 = (|$signed({(&{reg972})}));
              reg972 <= reg974[(4'hd):(3'h4)];
              reg973 <= ($unsigned((~|$unsigned(wire963))) + ((~&reg978[(3'h6):(3'h4)]) ?
                  $unsigned($unsigned(reg973)) : $signed((((8'ha1) ?
                      (8'ha2) : reg977) > $signed(reg978)))));
              reg976 = {(~$signed(($unsigned(wire964) ?
                      reg973[(3'h4):(1'h0)] : (reg967 ? reg970 : reg968)))),
                  {(reg975 - reg975[(3'h4):(1'h0)])}};
            end
          if ($unsigned($unsigned((~^reg972))))
            begin
              reg978 = $unsigned({((reg973 ?
                      forvar969[(3'h5):(1'h0)] : (&forvar976)) < forvar969)});
              reg980 = (forvar976[(1'h0):(1'h0)] || (!(~|(reg969[(2'h2):(2'h2)] - (reg978 ?
                  reg975 : reg967)))));
              reg981 <= $signed(wire965[(1'h0):(1'h0)]);
            end
          else
            begin
              reg977 <= wire966[(4'h8):(3'h6)];
              reg978 = (8'hb8);
              reg979 <= (~^reg974[(2'h3):(2'h2)]);
            end
        end
    end
  always
    @(posedge clk) begin
      reg982 = ((-reg973) ~^ reg972[(3'h6):(1'h0)]);
      if ((+$unsigned(($unsigned((~|reg973)) ?
          reg972 : wire965[(2'h2):(2'h2)]))))
        begin
          for (forvar983 = (1'h0); (forvar983 < (2'h3)); forvar983 = (forvar983 + (1'h1)))
            begin
              reg984 = (reg977[(2'h3):(1'h0)] ?
                  ((~&((-(8'h9d)) ?
                          wire963[(4'ha):(2'h2)] : (reg979 ?
                              reg977 : (7'h47)))) ?
                      (-reg975[(1'h1):(1'h0)]) : (wire966[(2'h2):(1'h0)] ?
                          (~$unsigned(reg982)) : reg981)) : reg981);
              reg985 <= reg981;
              reg986 = (~&(^~wire965[(2'h2):(1'h0)]));
              reg987 = (reg986[(2'h3):(2'h3)] ?
                  {wire963[(1'h0):(1'h0)]} : {$unsigned($unsigned({forvar983}))});
              reg988 = {{(reg977[(1'h1):(1'h0)] ?
                          (^(reg985 ? reg972 : wire966)) : wire964),
                      $signed(reg987)},
                  $signed(reg970[(5'h15):(4'h8)])};
            end
        end
      else
        begin
          for (forvar983 = (1'h0); (forvar983 < (1'h0)); forvar983 = (forvar983 + (1'h1)))
            begin
              reg984 = (|reg970[(3'h7):(3'h5)]);
              reg986 = $unsigned((~|($unsigned(reg984) ?
                  (reg977[(1'h1):(1'h0)] ?
                      $signed((8'hbb)) : reg984) : reg986[(3'h4):(3'h4)])));
              reg989 <= (~^(-$signed(reg987)));
              reg990 = ({$signed($signed(reg988[(2'h2):(2'h2)]))} * (-reg974));
            end
          reg991 = $signed((+($unsigned({reg982}) ?
              reg970 : $signed((reg986 ? wire966 : reg974)))));
          reg992 <= {(((wire966[(4'hd):(2'h2)] ?
                  (reg985 ?
                      wire963 : reg987) : reg979[(1'h0):(1'h0)]) + (7'h48)) && (~$unsigned((reg970 - (8'had)))))};
        end
    end
  assign wire993 = reg992[(4'hc):(3'h6)];
  assign wire994 = ($unsigned($unsigned($unsigned(wire964[(4'h9):(3'h7)]))) >> $signed(wire963[(4'h9):(2'h2)]));
  assign wire995 = $signed(((reg981[(3'h6):(3'h5)] ?
                           (reg974 ?
                               $signed((8'hbd)) : (^reg975)) : $unsigned($signed(reg975))) ?
                       $signed(($unsigned(reg975) ?
                           (reg973 >> (8'ha3)) : (wire964 > reg981))) : $signed((+reg985))));
  assign wire996 = (+(~$unsigned(wire965)));
  always
    @(posedge clk) begin
      if ($signed($unsigned(($unsigned(wire993) >> $unsigned(reg973)))))
        begin
          reg997 <= (~((($signed(reg977) + wire964[(4'h9):(1'h0)]) ?
                  (wire994[(3'h5):(3'h5)] || {wire963,
                      (8'h9f)}) : (~|$unsigned(reg977))) ?
              reg970[(4'ha):(4'h8)] : {(wire964 == (wire994 ?
                      wire964 : (8'h9d)))}));
          for (forvar998 = (1'h0); (forvar998 < (1'h1)); forvar998 = (forvar998 + (1'h1)))
            begin
              reg999 <= (^wire964);
              reg1000 = $signed($signed({reg997}));
              reg1001 = (reg974[(1'h0):(1'h0)] ?
                  (+forvar998[(4'he):(3'h6)]) : reg975);
            end
          for (forvar1002 = (1'h0); (forvar1002 < (1'h0)); forvar1002 = (forvar1002 + (1'h1)))
            begin
              reg1003 = reg975[(1'h0):(1'h0)];
              reg1004 <= (&($unsigned({reg975[(2'h2):(2'h2)]}) & forvar998[(3'h4):(1'h0)]));
              reg1005 <= reg997[(2'h2):(1'h0)];
              reg1006 = $unsigned($unsigned($unsigned(((reg970 && wire964) ^~ reg977))));
            end
          reg1007 <= $unsigned((((wire964 ?
              {wire995} : (forvar998 + (8'hbb))) & ($signed(reg970) & $unsigned(reg992))) + $unsigned(wire995[(1'h1):(1'h0)])));
          if (reg973)
            begin
              reg1008 = {((((~reg1004) + wire995[(1'h1):(1'h1)]) ?
                          reg1004 : ({reg1005} ?
                              reg1000 : $signed(forvar1002))) ?
                      (reg1007[(3'h4):(1'h1)] <= (|$unsigned(reg1007))) : wire996[(2'h3):(1'h0)])};
            end
          else
            begin
              reg1009 <= ((-$signed(wire966)) << ($unsigned(($unsigned(forvar1002) >= reg1006)) ?
                  (^$unsigned({(7'h42)})) : reg977));
              reg1010 <= reg974[(1'h1):(1'h0)];
            end
        end
      else
        begin
          for (forvar997 = (1'h0); (forvar997 < (1'h1)); forvar997 = (forvar997 + (1'h1)))
            begin
              reg998 <= (~$unsigned((($signed(reg975) ?
                  (~&forvar998) : $signed(reg1004)) >>> reg1003[(2'h2):(2'h2)])));
              reg999 <= ($signed((($signed(reg1010) ? reg1007 : reg1000) ?
                      reg979 : $signed(reg974[(2'h3):(2'h3)]))) ?
                  {(^~reg977[(1'h1):(1'h0)])} : $signed(wire993));
              reg1002 <= $signed((-(wire965[(1'h1):(1'h0)] ?
                  (reg997[(4'hd):(4'h8)] ?
                      {(8'ha9)} : $unsigned(reg973)) : (|$signed(reg975)))));
              reg1004 <= {reg970[(5'h16):(5'h13)]};
              reg1005 <= reg1003[(1'h0):(1'h0)];
            end
        end
      for (forvar1011 = (1'h0); (forvar1011 < (1'h1)); forvar1011 = (forvar1011 + (1'h1)))
        begin
          if (forvar1002)
            begin
              reg1012 <= (((reg977[(1'h1):(1'h0)] || {(|reg985)}) ?
                  $unsigned(reg1010[(3'h7):(1'h0)]) : ($unsigned(reg1008[(1'h1):(1'h1)]) != (!{reg1007}))) <= (((wire966 * $signed((8'hbe))) ?
                  (+(reg1004 ?
                      forvar1011 : (8'h9d))) : (-reg1002[(1'h1):(1'h0)])) <= (reg997 ?
                  ($unsigned(wire994) != reg970[(4'ha):(1'h0)]) : $signed(forvar1002[(4'ha):(3'h4)]))));
              reg1013 <= {(wire966 ^~ $unsigned($unsigned(reg1005)))};
            end
          else
            begin
              reg1014 = (~^wire965[(2'h2):(1'h1)]);
              reg1015 <= ((($unsigned($unsigned(forvar1011)) ?
                      $signed(wire964[(4'hb):(3'h5)]) : (|(~^reg972))) >= {{reg973[(3'h7):(3'h4)],
                          (wire964 ? reg985 : reg1012)},
                      $signed($signed(forvar997))}) ?
                  $signed((((reg975 ?
                          reg981 : reg1012) <<< (wire993 && wire994)) ?
                      forvar997[(5'h13):(4'hf)] : (~|reg1007))) : (~reg1012));
              reg1016 <= reg1004[(1'h0):(1'h0)];
            end
          reg1017 = $unsigned(reg1004);
        end
      reg1018 = ({(8'ha2)} ? wire996 : $unsigned($unsigned((+(~|reg972)))));
    end
  always
    @(posedge clk) begin
      if (reg979)
        begin
          reg1019 = {$signed(reg1009[(1'h1):(1'h0)])};
        end
      else
        begin
          reg1019 = ($unsigned((-wire966[(3'h7):(3'h6)])) ~^ (~^(^~($signed(wire993) >= reg974))));
          if ((({(^reg974[(4'hc):(2'h3)]), ($unsigned((8'hb6)) >> (+(8'hb2)))} ?
                  $signed((!$signed((7'h48)))) : $signed((~^reg1019[(5'h10):(2'h2)]))) ?
              (~^$unsigned($signed($unsigned((8'hac))))) : (|reg989)))
            begin
              reg1020 <= $unsigned((reg970 ?
                  (wire996 | $signed((reg1012 ?
                      reg974 : reg1019))) : reg975[(2'h2):(1'h0)]));
              reg1021 <= reg975;
              reg1022 = (reg970[(3'h5):(3'h4)] ?
                  reg997[(4'hb):(4'h9)] : reg992[(3'h7):(3'h7)]);
            end
          else
            begin
              reg1022 = (+reg974);
              reg1023 = ($signed((-(((8'hb4) ?
                  reg981 : wire965) * (wire963 && (8'ha1))))) <= $signed(reg973));
              reg1024 <= (^((8'ha6) + $unsigned((~^reg977[(1'h1):(1'h0)]))));
              reg1025 = ($unsigned((8'hac)) ?
                  (!({$signed(reg1024),
                      (+wire965)} ~^ reg970[(3'h6):(3'h5)])) : reg1013[(1'h0):(1'h0)]);
            end
          if ((((((&reg999) ? (reg1015 ? reg1010 : (8'hb5)) : (7'h43)) ?
                  reg1015[(4'hb):(4'ha)] : ($unsigned(reg1022) ?
                      $unsigned(reg1009) : $signed(wire965))) ?
              (^(~&$signed(reg1021))) : (((~|wire964) ?
                      (reg1002 < reg1016) : (wire995 >= reg1007)) ?
                  $unsigned(((8'hb3) ?
                      wire993 : reg970)) : $signed(reg1002))) >> (~(|(8'hb6)))))
            begin
              reg1026 <= $signed($unsigned((($signed(wire966) ~^ wire965) ?
                  $unsigned((reg977 << (7'h41))) : ((wire996 ?
                      wire994 : (8'hb0)) ^ reg975[(1'h1):(1'h0)]))));
              reg1027 = wire963;
              reg1028 <= reg1012[(2'h2):(1'h1)];
              reg1029 = (((8'hb0) == reg1023) ?
                  $signed({$unsigned((reg1022 ?
                          (8'hbd) : reg1027))}) : $unsigned($signed(($unsigned(reg1016) ?
                      $signed(reg998) : ((8'hb5) ? reg975 : wire994)))));
            end
          else
            begin
              reg1027 = ((+$unsigned($unsigned(reg997))) >> (8'ha9));
              reg1029 = (wire995 < reg1016);
              reg1030 <= (reg970[(3'h7):(2'h2)] || ((((8'h9f) ^~ reg1005) ?
                  {reg977, (+reg972)} : reg1007) - wire965[(2'h2):(2'h2)]));
              reg1031 = $unsigned(((($signed(wire994) ?
                      reg999[(3'h5):(2'h2)] : reg972[(4'h8):(3'h4)]) - ($unsigned((7'h4a)) ?
                      (!wire993) : (-reg992))) ?
                  $signed(({reg989} != $signed(reg989))) : (((|(8'ha2)) ?
                          $unsigned(reg1010) : $signed(reg1025)) ?
                      $unsigned($signed(reg999)) : reg1012)));
            end
          if ($unsigned($signed($signed({$unsigned(reg998)}))))
            begin
              reg1032 = {$signed(((-(~|reg992)) >> (|wire993)))};
              reg1033 <= wire966;
              reg1034 = $signed(wire996[(2'h2):(1'h0)]);
            end
          else
            begin
              reg1033 <= (8'ha0);
              reg1034 = (reg998[(3'h4):(2'h3)] <= reg974);
              reg1035 <= ({$unsigned({reg1032, reg973[(3'h4):(1'h0)]})} ?
                  $signed((wire965 ?
                      (reg1032 <<< (wire966 < reg1032)) : $unsigned((reg1004 <<< wire995)))) : $unsigned($signed($signed((!reg1020)))));
              reg1036 <= reg1024;
            end
          reg1037 <= (reg1033 ?
              ({(+reg1002[(3'h4):(2'h3)])} ?
                  reg1025 : ($signed((reg1016 ^~ reg970)) >> {reg1021,
                      reg998[(1'h1):(1'h0)]})) : ((({wire993} ?
                      $signed((8'ha7)) : (reg981 >>> reg975)) ?
                  reg1013[(1'h1):(1'h1)] : (&(reg1030 ?
                      reg1036 : reg1013))) || reg1032));
        end
      reg1038 <= reg992;
      if ((reg989 ^~ reg1024))
        begin
          reg1039 = ((8'h9d) >= ($signed($unsigned({reg1004})) & $signed({reg1019[(5'h17):(3'h7)]})));
          for (forvar1040 = (1'h0); (forvar1040 < (2'h3)); forvar1040 = (forvar1040 + (1'h1)))
            begin
              reg1041 = ((reg1027[(1'h0):(1'h0)] ?
                  ($signed({forvar1040}) ?
                      $signed($unsigned(reg1037)) : {(^(8'hb7)),
                          (reg1010 ?
                              reg1034 : reg1005)}) : (~&reg998)) >>> {reg1020,
                  wire993});
            end
          if (($unsigned((+(reg1034 || $unsigned((8'ha5))))) ?
              ($signed(((reg1025 ?
                  reg1020 : reg1010) <<< (~^reg1004))) >>> $signed(reg1015)) : (~^reg1026[(3'h6):(2'h2)])))
            begin
              reg1042 <= reg1025[(3'h5):(1'h1)];
              reg1043 <= reg1041[(4'hc):(4'hb)];
              reg1044 = reg1038[(3'h7):(1'h1)];
            end
          else
            begin
              reg1042 <= reg1043[(1'h1):(1'h0)];
            end
          reg1045 <= (reg1029 | (!$unsigned($unsigned(reg1015[(3'h6):(2'h3)]))));
        end
      else
        begin
          reg1040 <= (reg998[(3'h6):(2'h2)] ^ $unsigned(reg1036[(3'h7):(2'h3)]));
          for (forvar1041 = (1'h0); (forvar1041 < (2'h3)); forvar1041 = (forvar1041 + (1'h1)))
            begin
              reg1044 = $unsigned(reg1038[(3'h4):(1'h0)]);
              reg1045 <= (($unsigned($unsigned($signed(reg998))) ?
                  ($signed((wire963 + reg1033)) > (|reg1015)) : reg1041) != (&reg1042));
            end
          reg1046 = $signed(reg1015);
        end
    end
  always
    @(posedge clk) begin
      reg1047 = (-((reg1002[(1'h0):(1'h0)] > $signed(wire963)) ?
          reg1028 : $signed(reg1038[(3'h5):(1'h1)])));
      if ((~|wire965[(1'h0):(1'h0)]))
        begin
          reg1048 <= (reg1043[(3'h5):(1'h0)] ?
              $unsigned(reg979[(3'h6):(3'h4)]) : ((reg970[(4'hc):(4'ha)] ?
                      ($signed(wire996) ?
                          (reg1038 + reg1030) : {reg1005}) : $signed((reg989 ?
                          (7'h43) : (8'ha6)))) ?
                  ((8'h9c) <<< (~^$signed((8'ha4)))) : $unsigned(reg1037)));
        end
      else
        begin
          for (forvar1048 = (1'h0); (forvar1048 < (2'h2)); forvar1048 = (forvar1048 + (1'h1)))
            begin
              reg1049 = (((~(|(~reg1007))) ?
                  $signed({$unsigned((8'hbf)),
                      (reg1005 << reg1037)}) : reg992) > ((reg1033 && {wire963,
                      reg1021[(3'h4):(1'h1)]}) ?
                  ((^~(reg977 > (8'hba))) ^ ($unsigned((8'ha8)) ?
                      (-reg998) : reg972[(4'h8):(1'h0)])) : $signed({$signed(wire963)})));
              reg1050 <= wire996;
              reg1051 = $signed($signed(((-(~reg1040)) ?
                  reg1004[(2'h2):(1'h1)] : ((~&wire993) ?
                      $signed((8'hbc)) : reg970[(4'hc):(4'hc)]))));
              reg1052 = wire993[(4'h8):(2'h3)];
              reg1053 <= ({wire994[(2'h3):(1'h0)]} + (^~(8'ha8)));
            end
          for (forvar1054 = (1'h0); (forvar1054 < (2'h3)); forvar1054 = (forvar1054 + (1'h1)))
            begin
              reg1055 <= (^$signed((reg1048 <= reg1033[(4'h9):(4'h8)])));
            end
        end
    end
  assign wire1056 = (8'hb4);
  always
    @(posedge clk) begin
      if ($signed((reg1021[(3'h4):(2'h2)] << {({reg974, wire996} ^~ (wire965 ?
              reg999 : reg1036))})))
        begin
          for (forvar1057 = (1'h0); (forvar1057 < (2'h2)); forvar1057 = (forvar1057 + (1'h1)))
            begin
              reg1058 = ($unsigned(wire996) ?
                  ((7'h42) ?
                      wire994[(3'h5):(1'h1)] : (8'hb3)) : $unsigned($unsigned(($unsigned(reg997) >= ((8'hac) ?
                      reg1053 : reg985)))));
              reg1059 = (~|$unsigned((7'h41)));
              reg1060 = reg992;
              reg1061 = $unsigned($unsigned({$unsigned(reg973[(3'h7):(2'h3)]),
                  {reg1005[(3'h7):(3'h7)]}}));
              reg1062 = (($unsigned((~&(~reg981))) ?
                  reg1024[(3'h7):(2'h2)] : $unsigned(((~reg1036) ?
                      reg992 : reg1004))) >= (reg974[(4'h8):(2'h3)] ?
                  reg1061[(2'h3):(2'h2)] : (reg1020[(1'h0):(1'h0)] ?
                      $signed((reg1016 ?
                          wire963 : reg975)) : $signed($signed(reg1020)))));
            end
          if (((-(reg1045[(2'h3):(2'h2)] ^ (^~(!wire994)))) ?
              reg1028 : $unsigned(($unsigned($signed(wire993)) ?
                  reg1007 : (~|{reg1009, reg1036})))))
            begin
              reg1063 = $unsigned((~|$unsigned(((wire994 ?
                  (8'ha8) : reg970) ^~ (wire994 ? reg1016 : reg989)))));
              reg1064 = $signed($signed(reg977));
            end
          else
            begin
              reg1063 = {(^~(^(reg1059 ? $signed(reg1050) : reg1059))),
                  ((^~reg1010[(4'h8):(2'h2)]) ? (~&reg1033) : {(+(~(8'hb8)))})};
            end
          reg1065 = $signed((8'hb2));
          for (forvar1066 = (1'h0); (forvar1066 < (2'h2)); forvar1066 = (forvar1066 + (1'h1)))
            begin
              reg1067 <= {reg1045[(4'h9):(3'h5)]};
            end
        end
      else
        begin
          reg1057 = (-$signed((reg999[(1'h1):(1'h0)] && (~&reg1028))));
        end
      reg1068 = (((reg1028 ?
          reg972 : reg1060[(4'h9):(4'h9)]) | {(reg1020[(5'h17):(5'h17)] ?
              (reg999 >= reg979) : $unsigned(reg985))}) || reg974[(3'h7):(1'h0)]);
    end
  always
    @(posedge clk) begin
      if ($unsigned(reg1005[(3'h5):(1'h0)]))
        begin
          reg1069 = reg1040[(1'h1):(1'h1)];
          reg1070 <= $signed(reg974);
          for (forvar1071 = (1'h0); (forvar1071 < (2'h2)); forvar1071 = (forvar1071 + (1'h1)))
            begin
              reg1072 <= $signed($unsigned($signed(reg974[(4'hd):(4'hd)])));
              reg1073 <= $signed({reg1028[(3'h4):(3'h4)],
                  $unsigned(((-(8'hae)) ?
                      (reg1055 ? reg1012 : reg1055) : (reg985 ~^ reg1069)))});
              reg1074 <= {(-($signed(reg1038[(4'hc):(4'h9)]) ?
                      $unsigned(wire993[(5'h15):(4'hd)]) : reg1037[(2'h2):(1'h1)]))};
              reg1075 <= {reg1053};
            end
          reg1076 = {(^~reg1043),
              (!$signed({wire964, wire963[(1'h1):(1'h1)]}))};
        end
      else
        begin
          reg1070 <= (7'h49);
          reg1071 = reg1037[(4'hd):(3'h4)];
          if ($signed($unsigned($unsigned($unsigned((wire994 <= reg1043))))))
            begin
              reg1072 <= $unsigned({($unsigned(((8'hb4) & (7'h43))) + $unsigned($signed(reg1010)))});
              reg1073 <= $signed(reg1074);
            end
          else
            begin
              reg1076 = (|$signed($signed(reg1076[(3'h5):(3'h4)])));
              reg1077 = (($signed(reg1009) ?
                  $unsigned($signed(reg1024)) : $unsigned(reg997[(4'hc):(2'h2)])) ^ (reg1009 ?
                  (~^$unsigned($unsigned(wire964))) : reg1020));
              reg1078 <= (!reg1077[(4'h8):(2'h3)]);
              reg1079 = ((reg975[(1'h1):(1'h1)] - $signed(({reg1020, (8'hbe)} ?
                  (8'ha5) : $unsigned(reg1009)))) <<< reg1024);
              reg1080 <= $signed(((((reg1053 ? reg1028 : reg1015) ?
                  reg1043[(3'h4):(2'h3)] : wire966[(2'h2):(2'h2)]) + $signed(wire995[(4'h8):(3'h7)])) + {$signed((reg1067 ?
                      reg1071 : wire995)),
                  reg1076[(4'he):(1'h0)]}));
            end
          if (({$unsigned($unsigned((!(8'ha7)))),
              reg1069} <= (~^$signed(reg1078))))
            begin
              reg1081 = {((~^((reg1074 && reg998) ^ {reg1077})) ?
                      (+reg1013[(1'h1):(1'h0)]) : (((!reg972) >= reg1043) ?
                          $signed((~reg1043)) : $unsigned(((8'ha0) ^~ (8'hac)))))};
            end
          else
            begin
              reg1082 <= ($signed(reg1010) ?
                  (~|($signed($unsigned(reg970)) ?
                      reg1043 : (&$signed((8'hbb))))) : (reg1015 ?
                      reg1080[(1'h0):(1'h0)] : (-reg1002)));
            end
          for (forvar1083 = (1'h0); (forvar1083 < (3'h4)); forvar1083 = (forvar1083 + (1'h1)))
            begin
              reg1084 <= $unsigned(($signed($signed($signed(reg1080))) == wire965[(1'h0):(1'h0)]));
              reg1085 <= (reg1036[(3'h7):(3'h7)] ?
                  (((|reg1020[(5'h15):(3'h7)]) >>> (8'haa)) ?
                      reg1080 : ($unsigned((8'hab)) > ((reg1045 >>> (7'h45)) & ((8'ha8) ?
                          reg1030 : reg1071)))) : (reg1080 < (&({reg975,
                          wire1056} ?
                      (reg1026 ? reg1026 : reg1071) : reg974))));
              reg1086 = wire964;
            end
        end
      reg1087 <= (^~(8'ha0));
      reg1088 <= wire965;
      if (reg1050)
        begin
          if ($signed((8'ha6)))
            begin
              reg1089 = {{(|$unsigned(reg1079))}};
              reg1090 <= (8'hba);
            end
          else
            begin
              reg1089 = reg1028;
              reg1090 <= $unsigned({$unsigned($unsigned(((8'hab) * reg977)))});
              reg1091 <= reg977;
            end
        end
      else
        begin
          reg1090 <= reg970[(4'hb):(3'h6)];
          reg1091 <= (&forvar1083);
          for (forvar1092 = (1'h0); (forvar1092 < (1'h1)); forvar1092 = (forvar1092 + (1'h1)))
            begin
              reg1093 <= $unsigned($signed(((8'ha3) ?
                  (wire1056[(3'h6):(2'h3)] ?
                      reg973 : wire1056[(4'h8):(2'h2)]) : forvar1092)));
              reg1094 = ({({(|(8'hab))} ?
                      reg1038[(4'ha):(3'h4)] : reg1082[(4'h8):(4'h8)])} ~^ ($unsigned((+$unsigned(reg1040))) ?
                  $signed(reg1055) : reg1077[(5'h11):(4'hd)]));
              reg1095 = reg1026;
              reg1096 = (7'h48);
            end
          if ((($signed(reg1078) ?
                  reg1090[(2'h2):(1'h0)] : {$signed($signed(reg972))}) ?
              (~^wire966) : (wire966 == reg1053[(3'h4):(1'h0)])))
            begin
              reg1097 = {$signed(wire963),
                  ((((reg1040 ?
                          reg1020 : reg1002) <<< reg1028) << (reg1040[(1'h1):(1'h1)] >>> ((8'ha9) <= reg1082))) ?
                      reg1089[(3'h5):(1'h1)] : $signed({reg972[(3'h4):(1'h0)]}))};
              reg1098 = {((wire1056[(2'h2):(1'h1)] || {reg1067[(3'h5):(1'h1)]}) ?
                      $unsigned($signed((+wire994))) : $signed(reg1036[(3'h6):(2'h3)]))};
            end
          else
            begin
              reg1099 <= (&$unsigned(((~|(~reg1070)) ?
                  ($unsigned(reg975) ?
                      $signed((8'haf)) : $unsigned((7'h45))) : reg1013)));
              reg1100 = ({($unsigned((reg1035 - reg1067)) ?
                          reg1021[(1'h1):(1'h1)] : $signed({(8'ha9),
                              reg1004}))} ?
                  ((reg1033[(4'ha):(4'h9)] ?
                      $unsigned(forvar1071[(5'h10):(4'hb)]) : (8'hb3)) >> (reg970 ^ (~|(reg1088 || (8'hb3))))) : (({(~|reg1053),
                              (-reg1098)} ?
                          $unsigned((reg1085 ^~ reg1007)) : reg1033) ?
                      $unsigned({(reg1070 ?
                              reg1009 : reg1070)}) : reg1020[(5'h12):(1'h1)]));
              reg1101 = reg1082[(4'hf):(4'ha)];
              reg1102 = $signed($unsigned($unsigned((!reg1040))));
            end
        end
    end
  assign wire1103 = $unsigned({((wire964[(3'h5):(2'h2)] ?
                                $signed(reg1026) : (reg970 ?
                                    reg1090 : (8'hb7))) ?
                            $unsigned((wire965 ?
                                reg1080 : reg1091)) : ($signed(reg1026) ?
                                (reg979 ?
                                    reg1020 : reg1099) : wire965[(2'h2):(1'h1)]))});
  always
    @(posedge clk) begin
      reg1104 = (~$unsigned($unsigned({(~reg1033)})));
      if (((&({reg1004[(1'h0):(1'h0)],
          $signed(reg1090)} ~^ reg1072[(3'h6):(3'h6)])) != wire964))
        begin
          reg1105 <= $unsigned((^($signed({(7'h40),
              reg1021}) != (~&{(7'h41)}))));
          for (forvar1106 = (1'h0); (forvar1106 < (3'h4)); forvar1106 = (forvar1106 + (1'h1)))
            begin
              reg1107 = (8'ha6);
            end
        end
      else
        begin
          for (forvar1105 = (1'h0); (forvar1105 < (3'h4)); forvar1105 = (forvar1105 + (1'h1)))
            begin
              reg1106 = reg1070[(1'h0):(1'h0)];
            end
          reg1108 <= $unsigned(reg1009);
          if (wire964[(3'h7):(3'h4)])
            begin
              reg1109 <= (^~reg977);
              reg1110 = (8'h9e);
              reg1111 <= reg1055;
              reg1112 <= (~reg989);
              reg1113 <= $signed({((forvar1106 ?
                          ((8'hba) ? reg1050 : (8'hac)) : $unsigned(reg1015)) ?
                      $unsigned((reg1045 + reg972)) : ({(8'hbb),
                          reg1010} ^~ $signed(reg1042))),
                  (((reg1091 ? wire964 : (7'h4a)) >> (reg1070 ?
                      reg1038 : reg999)) & {(reg1040 ? reg977 : reg1045)})});
            end
          else
            begin
              reg1109 <= reg1112;
              reg1110 = $unsigned((~reg970));
              reg1114 = (reg1020[(5'h11):(5'h11)] ?
                  (+{$signed(reg1107[(2'h2):(1'h0)]),
                      $signed(((8'had) ?
                          reg1013 : reg1048))}) : (-{forvar1106}));
            end
          for (forvar1115 = (1'h0); (forvar1115 < (1'h0)); forvar1115 = (forvar1115 + (1'h1)))
            begin
              reg1116 <= (~^(8'ha2));
              reg1117 <= $signed(((wire1103 >= (reg979[(3'h4):(1'h1)] <<< reg974[(4'h8):(3'h6)])) != wire1103));
              reg1118 <= (&(^~reg1048[(3'h4):(1'h1)]));
              reg1119 <= reg1088[(4'hd):(4'h9)];
            end
          reg1120 <= (reg970 ?
              ($signed({wire966}) ?
                  reg1073[(3'h4):(2'h3)] : $signed(($unsigned(reg973) ?
                      (reg1035 + (8'hb4)) : (&reg1048)))) : (|reg1007));
        end
      reg1121 = (($unsigned(((~&reg1002) ? reg1043 : $signed(reg1009))) ?
              ($signed(reg1002[(2'h2):(1'h0)]) <= $unsigned((+(7'h49)))) : $unsigned((reg1118[(1'h0):(1'h0)] ?
                  (!(7'h42)) : (wire1103 ? reg1119 : reg1120)))) ?
          (reg1012 - reg1085) : ({reg1119, wire996} ?
              (wire963[(3'h5):(1'h1)] == reg1070) : reg979));
    end
  assign wire1122 = wire995;
  always
    @(posedge clk) begin
      reg1123 = (8'hbf);
      if ($signed((8'ha5)))
        begin
          reg1124 <= ((($unsigned((reg1075 || reg1070)) * (wire966 ?
                  {reg1091, wire1056} : reg992)) ?
              $unsigned(reg1112) : ($unsigned($signed(reg979)) << $signed((reg1112 & reg1085)))) != ((wire1056 <<< (reg981[(3'h7):(3'h6)] ?
                  ((8'hb6) ? reg1013 : reg1119) : $signed(wire1056))) ?
              $signed($unsigned((reg1070 & reg1078))) : ($unsigned($signed(wire965)) == reg1036)));
          reg1125 <= reg1087;
          reg1126 <= (((~|reg998) | (~&reg1117[(3'h5):(3'h5)])) << $unsigned($unsigned($unsigned((-reg1124)))));
          reg1127 <= $signed($signed({$signed(reg1005), reg1123}));
        end
      else
        begin
          reg1128 = (8'hbb);
          reg1129 = $unsigned((^~$signed((^~(reg989 ? reg1127 : reg1028)))));
          reg1130 = $signed($unsigned({(~^((8'had) >> (8'ha1))),
              ((!reg1082) ^~ {reg1080})}));
          for (forvar1131 = (1'h0); (forvar1131 < (3'h4)); forvar1131 = (forvar1131 + (1'h1)))
            begin
              reg1132 <= (^$unsigned(($unsigned($signed(reg1088)) ?
                  ({wire965} <<< $signed(reg1045)) : $unsigned(((7'h46) * wire996)))));
              reg1133 = wire1056[(2'h3):(2'h3)];
              reg1134 = reg1111[(5'h13):(3'h4)];
              reg1135 = reg1030;
              reg1136 = ((reg981[(3'h6):(3'h5)] ?
                      (reg1026[(1'h0):(1'h0)] <= $unsigned($signed(reg1105))) : (({(8'ha7),
                              reg1111} ?
                          reg1026[(4'h8):(1'h1)] : (reg1130 << reg972)) << (reg1007[(4'hf):(4'hd)] ?
                          $signed(reg1002) : wire996[(1'h1):(1'h0)]))) ?
                  $unsigned(reg1123[(4'h9):(1'h1)]) : (reg1091 || reg1012[(1'h1):(1'h1)]));
            end
          reg1137 = reg1132[(2'h2):(1'h1)];
        end
      reg1138 <= reg1005;
    end
  assign wire1139 = ((|{reg992}) && reg1002);
  assign wire1140 = ($signed((+reg1093)) & {$unsigned((~(reg1021 - wire965)))});
  assign wire1141 = $unsigned($unsigned((wire996[(3'h7):(2'h2)] ?
                        (~|((8'hb5) ?
                            reg1085 : reg1016)) : $signed((^~reg1075)))));
  assign wire1142 = wire993[(4'he):(4'hd)];
  always
    @(posedge clk) begin
      for (forvar1143 = (1'h0); (forvar1143 < (2'h2)); forvar1143 = (forvar1143 + (1'h1)))
        begin
          reg1144 = (!$signed($unsigned((-reg1111[(4'ha):(1'h0)]))));
        end
      reg1145 = (reg1118[(1'h0):(1'h0)] > (~|((8'haf) ?
          (-$unsigned(reg1072)) : (~&{reg1080}))));
      if ((reg1015[(5'h10):(4'h8)] ?
          {({((8'hb7) && reg1120),
                  reg1099[(2'h2):(2'h2)]} > ($signed(reg1084) >>> (reg989 ?
                  reg1048 : reg975))),
              {$signed(wire1056[(1'h0):(1'h0)]),
                  (reg970[(5'h15):(4'hf)] ?
                      {reg981} : (reg1004 >= reg1015))}} : ($signed(wire964) ?
              (^~{(reg1007 ?
                      reg1099 : reg1088)}) : ($unsigned((&reg1087)) + reg1040))))
        begin
          for (forvar1146 = (1'h0); (forvar1146 < (1'h0)); forvar1146 = (forvar1146 + (1'h1)))
            begin
              reg1147 <= reg1005;
              reg1148 = $signed({$unsigned(($signed(reg1013) ?
                      $signed((8'hbb)) : wire994[(2'h3):(2'h3)]))});
              reg1149 <= (!({$signed(reg1042),
                  {(reg1085 ? (7'h43) : (8'ha3)),
                      $signed((8'hb4))}} >= reg1148[(4'h8):(1'h0)]));
            end
          for (forvar1150 = (1'h0); (forvar1150 < (1'h1)); forvar1150 = (forvar1150 + (1'h1)))
            begin
              reg1151 = (8'ha2);
              reg1152 <= (+reg1053[(2'h2):(1'h0)]);
              reg1153 <= {{(!({reg1148, (8'hbc)} != (!reg1037))),
                      $signed((-reg1070))}};
              reg1154 = (reg970[(4'hc):(4'h8)] ?
                  reg1147[(4'ha):(1'h0)] : (($signed((~^reg1125)) ?
                          (~|(wire993 <<< reg1053)) : (~^((8'hbf) >>> (7'h45)))) ?
                      {({reg1127,
                              reg1120} ^ $unsigned(reg1007))} : $unsigned((8'haf))));
              reg1155 <= $signed((&({reg1073} | (~$signed(reg1090)))));
            end
          for (forvar1156 = (1'h0); (forvar1156 < (3'h4)); forvar1156 = (forvar1156 + (1'h1)))
            begin
              reg1157 <= reg1016[(4'h8):(1'h0)];
            end
        end
      else
        begin
          if ($unsigned(($signed({$unsigned(wire1139)}) + (^reg998))))
            begin
              reg1146 = ($unsigned($unsigned(reg1124)) ?
                  wire1056 : $signed($unsigned(reg1036[(3'h6):(3'h5)])));
              reg1148 = reg1132;
            end
          else
            begin
              reg1147 <= reg1155[(5'h17):(4'h9)];
              reg1148 = reg1030[(3'h7):(1'h1)];
            end
          for (forvar1149 = (1'h0); (forvar1149 < (1'h1)); forvar1149 = (forvar1149 + (1'h1)))
            begin
              reg1150 = reg1113[(1'h0):(1'h0)];
              reg1151 = $signed(reg1050[(3'h5):(3'h5)]);
              reg1154 = $unsigned((-(7'h40)));
              reg1156 = {{reg1042}, reg989[(4'hc):(4'h9)]};
            end
          for (forvar1157 = (1'h0); (forvar1157 < (1'h1)); forvar1157 = (forvar1157 + (1'h1)))
            begin
              reg1158 <= (8'h9c);
              reg1159 <= (reg1105[(3'h5):(3'h5)] << (!(reg1013[(2'h3):(1'h1)] ?
                  ((~&reg981) & reg1033) : ($unsigned(reg1072) << {reg981,
                      reg1127}))));
            end
          reg1160 = (reg1156 ?
              $signed(reg1125[(1'h1):(1'h1)]) : ($unsigned($signed((reg1155 ?
                      reg1015 : reg1050))) ?
                  (+(7'h48)) : (^~(reg1157[(3'h4):(1'h0)] | $unsigned(reg1148)))));
        end
      reg1161 <= reg1012[(2'h2):(1'h1)];
      reg1162 <= (8'ha0);
    end
endmodule

(* use_dsp48="no" *) (* use_dsp="no" *) module module643
#(parameter param959 = (~&((((!(8'hbd)) > ((8'hb1) << (8'hbb))) - (((8'h9d) >> (7'h41)) ? (~|(8'had)) : ((8'hbf) ? (8'h9f) : (8'hb5)))) ^~ (~^{(-(8'hb1))}))))
(y, clk, wire648, wire647, wire646, wire645, wire644);
  output wire [(32'h1150):(32'h0)] y;
  input wire [(1'h0):(1'h0)] clk;
  input wire signed [(5'h12):(1'h0)] wire648;
  input wire [(4'ha):(1'h0)] wire647;
  input wire signed [(3'h5):(1'h0)] wire646;
  input wire [(4'h9):(1'h0)] wire645;
  input wire signed [(3'h6):(1'h0)] wire644;
  wire [(4'ha):(1'h0)] wire958;
  wire signed [(5'h18):(1'h0)] wire930;
  wire signed [(4'hd):(1'h0)] wire870;
  wire signed [(3'h6):(1'h0)] wire845;
  wire [(5'h17):(1'h0)] wire844;
  wire signed [(4'h9):(1'h0)] wire700;
  wire signed [(4'hd):(1'h0)] wire699;
  wire [(4'h9):(1'h0)] wire698;
  wire [(5'h17):(1'h0)] wire652;
  wire [(4'ha):(1'h0)] wire649;
  reg [(4'he):(1'h0)] reg956 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg955 = (1'h0);
  reg [(5'h17):(1'h0)] reg954 = (1'h0);
  reg [(5'h10):(1'h0)] reg952 = (1'h0);
  reg [(3'h4):(1'h0)] reg948 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg942 = (1'h0);
  reg [(3'h4):(1'h0)] reg945 = (1'h0);
  reg [(3'h6):(1'h0)] reg943 = (1'h0);
  reg [(3'h5):(1'h0)] reg940 = (1'h0);
  reg [(4'he):(1'h0)] reg937 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg936 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg935 = (1'h0);
  reg [(3'h4):(1'h0)] reg933 = (1'h0);
  reg [(5'h15):(1'h0)] reg932 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg929 = (1'h0);
  reg [(3'h4):(1'h0)] reg928 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg927 = (1'h0);
  reg [(5'h14):(1'h0)] reg925 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg923 = (1'h0);
  reg signed [(4'he):(1'h0)] reg922 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg919 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg916 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg913 = (1'h0);
  reg [(5'h13):(1'h0)] reg912 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg909 = (1'h0);
  reg [(5'h14):(1'h0)] reg907 = (1'h0);
  reg [(4'hf):(1'h0)] reg902 = (1'h0);
  reg [(5'h16):(1'h0)] reg901 = (1'h0);
  reg [(4'hb):(1'h0)] reg900 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg898 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg895 = (1'h0);
  reg [(4'hb):(1'h0)] reg894 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg891 = (1'h0);
  reg [(5'h12):(1'h0)] reg889 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg887 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg879 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg876 = (1'h0);
  reg [(5'h13):(1'h0)] reg875 = (1'h0);
  reg [(5'h12):(1'h0)] reg873 = (1'h0);
  reg [(4'he):(1'h0)] reg871 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg869 = (1'h0);
  reg [(4'ha):(1'h0)] reg866 = (1'h0);
  reg [(2'h3):(1'h0)] reg857 = (1'h0);
  reg [(5'h15):(1'h0)] reg856 = (1'h0);
  reg signed [(4'he):(1'h0)] reg854 = (1'h0);
  reg [(5'h13):(1'h0)] reg853 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg849 = (1'h0);
  reg [(4'hd):(1'h0)] reg847 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg841 = (1'h0);
  reg [(3'h4):(1'h0)] reg839 = (1'h0);
  reg signed [(4'he):(1'h0)] reg820 = (1'h0);
  reg [(4'hd):(1'h0)] reg836 = (1'h0);
  reg [(4'ha):(1'h0)] reg833 = (1'h0);
  reg [(4'ha):(1'h0)] reg832 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg830 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg829 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg828 = (1'h0);
  reg [(4'he):(1'h0)] reg824 = (1'h0);
  reg [(5'h17):(1'h0)] reg822 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg821 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg817 = (1'h0);
  reg [(4'ha):(1'h0)] reg815 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg814 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg813 = (1'h0);
  reg [(5'h12):(1'h0)] reg812 = (1'h0);
  reg [(2'h3):(1'h0)] reg810 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg807 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg806 = (1'h0);
  reg [(5'h14):(1'h0)] reg805 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg804 = (1'h0);
  reg [(5'h17):(1'h0)] reg803 = (1'h0);
  reg [(3'h4):(1'h0)] reg800 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg785 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg794 = (1'h0);
  reg [(2'h2):(1'h0)] reg792 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg791 = (1'h0);
  reg [(4'hb):(1'h0)] reg790 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg789 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg788 = (1'h0);
  reg [(4'ha):(1'h0)] reg786 = (1'h0);
  reg [(3'h7):(1'h0)] reg784 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg779 = (1'h0);
  reg [(4'hd):(1'h0)] reg777 = (1'h0);
  reg [(2'h3):(1'h0)] reg772 = (1'h0);
  reg [(5'h13):(1'h0)] reg769 = (1'h0);
  reg [(5'h13):(1'h0)] reg768 = (1'h0);
  reg [(5'h11):(1'h0)] reg767 = (1'h0);
  reg [(5'h12):(1'h0)] reg765 = (1'h0);
  reg [(3'h6):(1'h0)] reg762 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg761 = (1'h0);
  reg [(4'hc):(1'h0)] reg760 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg758 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg757 = (1'h0);
  reg [(5'h14):(1'h0)] reg755 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg754 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg753 = (1'h0);
  reg [(3'h7):(1'h0)] reg752 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg743 = (1'h0);
  reg signed [(3'h6):(1'h0)] reg741 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg736 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg738 = (1'h0);
  reg [(4'h9):(1'h0)] reg737 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg728 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg726 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg725 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg719 = (1'h0);
  reg [(4'hf):(1'h0)] reg723 = (1'h0);
  reg [(4'hb):(1'h0)] reg722 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg720 = (1'h0);
  reg [(5'h17):(1'h0)] reg718 = (1'h0);
  reg [(5'h17):(1'h0)] reg716 = (1'h0);
  reg [(4'ha):(1'h0)] reg715 = (1'h0);
  reg [(4'hb):(1'h0)] reg714 = (1'h0);
  reg [(5'h15):(1'h0)] reg712 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg710 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg709 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg706 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg695 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg693 = (1'h0);
  reg [(4'h8):(1'h0)] reg691 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg685 = (1'h0);
  reg [(5'h18):(1'h0)] reg689 = (1'h0);
  reg [(3'h6):(1'h0)] reg687 = (1'h0);
  reg [(4'h8):(1'h0)] reg686 = (1'h0);
  reg signed [(2'h2):(1'h0)] reg682 = (1'h0);
  reg [(5'h15):(1'h0)] reg681 = (1'h0);
  reg [(4'h8):(1'h0)] reg678 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg676 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg675 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg670 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg669 = (1'h0);
  reg [(3'h4):(1'h0)] reg667 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg666 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg665 = (1'h0);
  reg [(5'h10):(1'h0)] reg663 = (1'h0);
  reg [(3'h7):(1'h0)] reg658 = (1'h0);
  reg [(3'h6):(1'h0)] reg657 = (1'h0);
  reg [(4'h8):(1'h0)] reg656 = (1'h0);
  reg [(4'hb):(1'h0)] reg654 = (1'h0);
  reg [(4'hc):(1'h0)] reg653 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg651 = (1'h0);
  reg [(4'h8):(1'h0)] reg957 = (1'h0);
  reg [(4'ha):(1'h0)] reg953 = (1'h0);
  reg [(3'h6):(1'h0)] reg951 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg950 = (1'h0);
  reg [(5'h16):(1'h0)] reg949 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg947 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg944 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar938 = (1'h0);
  reg [(3'h5):(1'h0)] reg946 = (1'h0);
  reg [(4'he):(1'h0)] forvar944 = (1'h0);
  reg [(5'h10):(1'h0)] forvar942 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg941 = (1'h0);
  reg [(3'h4):(1'h0)] reg939 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg938 = (1'h0);
  reg signed [(5'h11):(1'h0)] forvar934 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg931 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg926 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg924 = (1'h0);
  reg [(5'h11):(1'h0)] reg921 = (1'h0);
  reg [(4'hd):(1'h0)] reg920 = (1'h0);
  reg signed [(2'h2):(1'h0)] forvar918 = (1'h0);
  reg [(5'h10):(1'h0)] forvar911 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg910 = (1'h0);
  reg [(2'h2):(1'h0)] reg917 = (1'h0);
  reg [(3'h7):(1'h0)] reg915 = (1'h0);
  reg [(4'hd):(1'h0)] reg914 = (1'h0);
  reg [(3'h7):(1'h0)] reg911 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar910 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg908 = (1'h0);
  reg [(3'h5):(1'h0)] reg906 = (1'h0);
  reg [(2'h3):(1'h0)] forvar905 = (1'h0);
  reg [(4'he):(1'h0)] reg904 = (1'h0);
  reg [(4'hf):(1'h0)] reg903 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar899 = (1'h0);
  reg [(3'h4):(1'h0)] reg897 = (1'h0);
  reg [(4'ha):(1'h0)] reg896 = (1'h0);
  reg signed [(5'h14):(1'h0)] forvar893 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg892 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg890 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg888 = (1'h0);
  reg signed [(4'he):(1'h0)] reg886 = (1'h0);
  reg signed [(4'ha):(1'h0)] reg885 = (1'h0);
  reg [(4'he):(1'h0)] reg884 = (1'h0);
  reg [(5'h18):(1'h0)] reg883 = (1'h0);
  reg [(4'hc):(1'h0)] reg882 = (1'h0);
  reg [(5'h10):(1'h0)] forvar881 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg880 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar878 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg877 = (1'h0);
  reg [(5'h17):(1'h0)] reg874 = (1'h0);
  reg [(3'h4):(1'h0)] reg872 = (1'h0);
  reg signed [(5'h16):(1'h0)] reg868 = (1'h0);
  reg [(4'he):(1'h0)] reg867 = (1'h0);
  reg signed [(5'h12):(1'h0)] reg865 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg864 = (1'h0);
  reg [(3'h5):(1'h0)] reg863 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar862 = (1'h0);
  reg [(5'h11):(1'h0)] reg861 = (1'h0);
  reg [(5'h14):(1'h0)] forvar860 = (1'h0);
  reg signed [(4'h8):(1'h0)] reg859 = (1'h0);
  reg signed [(5'h15):(1'h0)] reg848 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg858 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg855 = (1'h0);
  reg [(4'hb):(1'h0)] reg852 = (1'h0);
  reg [(2'h3):(1'h0)] reg851 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg850 = (1'h0);
  reg signed [(4'hb):(1'h0)] forvar848 = (1'h0);
  reg [(5'h18):(1'h0)] reg846 = (1'h0);
  reg [(4'h8):(1'h0)] reg843 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg842 = (1'h0);
  reg [(5'h14):(1'h0)] reg840 = (1'h0);
  reg signed [(5'h17):(1'h0)] forvar838 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar837 = (1'h0);
  reg [(5'h13):(1'h0)] reg825 = (1'h0);
  reg [(5'h11):(1'h0)] forvar821 = (1'h0);
  reg [(4'hf):(1'h0)] reg835 = (1'h0);
  reg [(5'h11):(1'h0)] reg834 = (1'h0);
  reg signed [(4'ha):(1'h0)] forvar831 = (1'h0);
  reg signed [(4'hc):(1'h0)] reg827 = (1'h0);
  reg [(4'he):(1'h0)] reg826 = (1'h0);
  reg signed [(4'h9):(1'h0)] forvar825 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg823 = (1'h0);
  reg [(4'he):(1'h0)] forvar820 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg819 = (1'h0);
  reg [(3'h6):(1'h0)] reg818 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg816 = (1'h0);
  reg [(5'h13):(1'h0)] reg811 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar809 = (1'h0);
  reg [(4'hc):(1'h0)] forvar808 = (1'h0);
  reg [(3'h6):(1'h0)] reg802 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg801 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg799 = (1'h0);
  reg [(4'hb):(1'h0)] reg798 = (1'h0);
  reg [(5'h15):(1'h0)] reg797 = (1'h0);
  reg [(4'ha):(1'h0)] forvar796 = (1'h0);
  reg [(5'h18):(1'h0)] reg795 = (1'h0);
  reg [(4'hb):(1'h0)] reg793 = (1'h0);
  reg [(5'h13):(1'h0)] reg787 = (1'h0);
  reg signed [(3'h5):(1'h0)] forvar785 = (1'h0);
  reg [(3'h5):(1'h0)] reg783 = (1'h0);
  reg [(4'hb):(1'h0)] forvar782 = (1'h0);
  reg [(4'h8):(1'h0)] reg781 = (1'h0);
  reg signed [(5'h13):(1'h0)] reg780 = (1'h0);
  reg [(4'hc):(1'h0)] reg778 = (1'h0);
  reg [(5'h11):(1'h0)] forvar776 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg775 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg774 = (1'h0);
  reg [(5'h14):(1'h0)] reg773 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg771 = (1'h0);
  reg [(4'he):(1'h0)] forvar770 = (1'h0);
  reg signed [(3'h4):(1'h0)] reg766 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar764 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg763 = (1'h0);
  reg [(4'hd):(1'h0)] reg759 = (1'h0);
  reg signed [(5'h10):(1'h0)] forvar757 = (1'h0);
  reg [(5'h13):(1'h0)] reg756 = (1'h0);
  reg [(3'h7):(1'h0)] reg749 = (1'h0);
  reg [(2'h3):(1'h0)] forvar748 = (1'h0);
  reg [(2'h2):(1'h0)] reg751 = (1'h0);
  reg [(2'h2):(1'h0)] reg750 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar749 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg748 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg747 = (1'h0);
  reg [(4'he):(1'h0)] reg746 = (1'h0);
  reg signed [(4'hd):(1'h0)] forvar745 = (1'h0);
  reg signed [(4'hd):(1'h0)] reg744 = (1'h0);
  reg [(5'h16):(1'h0)] reg742 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg733 = (1'h0);
  reg [(3'h5):(1'h0)] reg740 = (1'h0);
  reg [(4'hc):(1'h0)] reg739 = (1'h0);
  reg signed [(3'h4):(1'h0)] forvar736 = (1'h0);
  reg [(5'h15):(1'h0)] reg735 = (1'h0);
  reg [(2'h3):(1'h0)] reg734 = (1'h0);
  reg [(3'h4):(1'h0)] forvar733 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg732 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar731 = (1'h0);
  reg signed [(5'h16):(1'h0)] forvar730 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg729 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg727 = (1'h0);
  reg [(3'h7):(1'h0)] reg724 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar720 = (1'h0);
  reg [(5'h13):(1'h0)] forvar718 = (1'h0);
  reg signed [(4'he):(1'h0)] reg717 = (1'h0);
  reg signed [(4'he):(1'h0)] reg721 = (1'h0);
  reg signed [(2'h3):(1'h0)] forvar719 = (1'h0);
  reg signed [(3'h6):(1'h0)] forvar717 = (1'h0);
  reg signed [(4'hb):(1'h0)] reg713 = (1'h0);
  reg signed [(4'h9):(1'h0)] reg711 = (1'h0);
  reg signed [(5'h17):(1'h0)] reg708 = (1'h0);
  reg [(5'h16):(1'h0)] reg707 = (1'h0);
  reg signed [(3'h7):(1'h0)] reg705 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg704 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg703 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg702 = (1'h0);
  reg [(4'hf):(1'h0)] reg701 = (1'h0);
  reg [(5'h14):(1'h0)] reg697 = (1'h0);
  reg [(4'h8):(1'h0)] reg696 = (1'h0);
  reg [(5'h10):(1'h0)] reg694 = (1'h0);
  reg signed [(2'h3):(1'h0)] reg692 = (1'h0);
  reg [(4'hb):(1'h0)] reg688 = (1'h0);
  reg [(2'h3):(1'h0)] reg683 = (1'h0);
  reg signed [(5'h14):(1'h0)] reg690 = (1'h0);
  reg [(3'h7):(1'h0)] forvar688 = (1'h0);
  reg signed [(4'he):(1'h0)] forvar685 = (1'h0);
  reg [(5'h10):(1'h0)] reg684 = (1'h0);
  reg signed [(5'h13):(1'h0)] forvar683 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg680 = (1'h0);
  reg [(3'h4):(1'h0)] reg679 = (1'h0);
  reg [(5'h10):(1'h0)] reg677 = (1'h0);
  reg [(4'hb):(1'h0)] reg674 = (1'h0);
  reg [(5'h15):(1'h0)] reg673 = (1'h0);
  reg signed [(5'h18):(1'h0)] forvar672 = (1'h0);
  reg signed [(3'h5):(1'h0)] reg671 = (1'h0);
  reg signed [(5'h11):(1'h0)] reg668 = (1'h0);
  reg [(3'h7):(1'h0)] reg664 = (1'h0);
  reg [(4'hf):(1'h0)] reg662 = (1'h0);
  reg [(5'h15):(1'h0)] reg661 = (1'h0);
  reg signed [(5'h10):(1'h0)] reg660 = (1'h0);
  reg [(5'h12):(1'h0)] reg659 = (1'h0);
  reg signed [(4'hf):(1'h0)] forvar653 = (1'h0);
  reg signed [(4'hf):(1'h0)] reg655 = (1'h0);
  reg signed [(5'h18):(1'h0)] reg650 = (1'h0);
  assign y = {wire958,
                 wire930,
                 wire870,
                 wire845,
                 wire844,
                 wire700,
                 wire699,
                 wire698,
                 wire652,
                 wire649,
                 reg956,
                 reg955,
                 reg954,
                 reg952,
                 reg948,
                 reg942,
                 reg945,
                 reg943,
                 reg940,
                 reg937,
                 reg936,
                 reg935,
                 reg933,
                 reg932,
                 reg929,
                 reg928,
                 reg927,
                 reg925,
                 reg923,
                 reg922,
                 reg919,
                 reg916,
                 reg913,
                 reg912,
                 reg909,
                 reg907,
                 reg902,
                 reg901,
                 reg900,
                 reg898,
                 reg895,
                 reg894,
                 reg891,
                 reg889,
                 reg887,
                 reg879,
                 reg876,
                 reg875,
                 reg873,
                 reg871,
                 reg869,
                 reg866,
                 reg857,
                 reg856,
                 reg854,
                 reg853,
                 reg849,
                 reg847,
                 reg841,
                 reg839,
                 reg820,
                 reg836,
                 reg833,
                 reg832,
                 reg830,
                 reg829,
                 reg828,
                 reg824,
                 reg822,
                 reg821,
                 reg817,
                 reg815,
                 reg814,
                 reg813,
                 reg812,
                 reg810,
                 reg807,
                 reg806,
                 reg805,
                 reg804,
                 reg803,
                 reg800,
                 reg785,
                 reg794,
                 reg792,
                 reg791,
                 reg790,
                 reg789,
                 reg788,
                 reg786,
                 reg784,
                 reg779,
                 reg777,
                 reg772,
                 reg769,
                 reg768,
                 reg767,
                 reg765,
                 reg762,
                 reg761,
                 reg760,
                 reg758,
                 reg757,
                 reg755,
                 reg754,
                 reg753,
                 reg752,
                 reg743,
                 reg741,
                 reg736,
                 reg738,
                 reg737,
                 reg728,
                 reg726,
                 reg725,
                 reg719,
                 reg723,
                 reg722,
                 reg720,
                 reg718,
                 reg716,
                 reg715,
                 reg714,
                 reg712,
                 reg710,
                 reg709,
                 reg706,
                 reg695,
                 reg693,
                 reg691,
                 reg685,
                 reg689,
                 reg687,
                 reg686,
                 reg682,
                 reg681,
                 reg678,
                 reg676,
                 reg675,
                 reg670,
                 reg669,
                 reg667,
                 reg666,
                 reg665,
                 reg663,
                 reg658,
                 reg657,
                 reg656,
                 reg654,
                 reg653,
                 reg651,
                 reg957,
                 reg953,
                 reg951,
                 reg950,
                 reg949,
                 reg947,
                 reg944,
                 forvar938,
                 reg946,
                 forvar944,
                 forvar942,
                 reg941,
                 reg939,
                 reg938,
                 forvar934,
                 reg931,
                 reg926,
                 reg924,
                 reg921,
                 reg920,
                 forvar918,
                 forvar911,
                 reg910,
                 reg917,
                 reg915,
                 reg914,
                 reg911,
                 forvar910,
                 reg908,
                 reg906,
                 forvar905,
                 reg904,
                 reg903,
                 forvar899,
                 reg897,
                 reg896,
                 forvar893,
                 reg892,
                 reg890,
                 reg888,
                 reg886,
                 reg885,
                 reg884,
                 reg883,
                 reg882,
                 forvar881,
                 reg880,
                 forvar878,
                 reg877,
                 reg874,
                 reg872,
                 reg868,
                 reg867,
                 reg865,
                 reg864,
                 reg863,
                 forvar862,
                 reg861,
                 forvar860,
                 reg859,
                 reg848,
                 reg858,
                 reg855,
                 reg852,
                 reg851,
                 reg850,
                 forvar848,
                 reg846,
                 reg843,
                 reg842,
                 reg840,
                 forvar838,
                 forvar837,
                 reg825,
                 forvar821,
                 reg835,
                 reg834,
                 forvar831,
                 reg827,
                 reg826,
                 forvar825,
                 reg823,
                 forvar820,
                 reg819,
                 reg818,
                 reg816,
                 reg811,
                 forvar809,
                 forvar808,
                 reg802,
                 reg801,
                 reg799,
                 reg798,
                 reg797,
                 forvar796,
                 reg795,
                 reg793,
                 reg787,
                 forvar785,
                 reg783,
                 forvar782,
                 reg781,
                 reg780,
                 reg778,
                 forvar776,
                 reg775,
                 reg774,
                 reg773,
                 reg771,
                 forvar770,
                 reg766,
                 forvar764,
                 reg763,
                 reg759,
                 forvar757,
                 reg756,
                 reg749,
                 forvar748,
                 reg751,
                 reg750,
                 forvar749,
                 reg748,
                 reg747,
                 reg746,
                 forvar745,
                 reg744,
                 reg742,
                 reg733,
                 reg740,
                 reg739,
                 forvar736,
                 reg735,
                 reg734,
                 forvar733,
                 reg732,
                 forvar731,
                 forvar730,
                 reg729,
                 reg727,
                 reg724,
                 forvar720,
                 forvar718,
                 reg717,
                 reg721,
                 forvar719,
                 forvar717,
                 reg713,
                 reg711,
                 reg708,
                 reg707,
                 reg705,
                 reg704,
                 reg703,
                 reg702,
                 reg701,
                 reg697,
                 reg696,
                 reg694,
                 reg692,
                 reg688,
                 reg683,
                 reg690,
                 forvar688,
                 forvar685,
                 reg684,
                 forvar683,
                 reg680,
                 reg679,
                 reg677,
                 reg674,
                 reg673,
                 forvar672,
                 reg671,
                 reg668,
                 reg664,
                 reg662,
                 reg661,
                 reg660,
                 reg659,
                 forvar653,
                 reg655,
                 reg650,
                 (1'h0)};
  assign wire649 = (+(~$signed($unsigned((wire645 ? (7'h47) : wire646)))));
  always
    @(posedge clk) begin
      reg650 = wire644[(3'h6):(1'h1)];
      reg651 <= {wire649[(3'h4):(1'h1)],
          {wire649,
              $unsigned((wire646[(2'h3):(2'h2)] ?
                  wire647 : $signed((8'ha0))))}};
    end
  assign wire652 = $unsigned((&(wire645 > $unsigned(reg651))));
  always
    @(posedge clk) begin
      if (wire646)
        begin
          reg653 <= (wire649 ~^ (8'ha7));
          reg654 <= (&{($signed(wire652) < wire652), wire646[(1'h0):(1'h0)]});
          reg655 = ($signed((wire652 + $unsigned((wire648 * wire646)))) & $signed(($signed($signed(wire649)) << wire649)));
          if (wire649)
            begin
              reg656 <= $unsigned(reg651);
            end
          else
            begin
              reg656 <= $signed(wire645);
              reg657 <= ((reg653[(3'h4):(1'h1)] ?
                      {reg656, $signed(reg656)} : wire647[(4'ha):(4'h8)]) ?
                  $signed(wire648) : wire645);
              reg658 <= $unsigned((+(wire647 != wire649[(4'ha):(3'h7)])));
            end
        end
      else
        begin
          for (forvar653 = (1'h0); (forvar653 < (2'h3)); forvar653 = (forvar653 + (1'h1)))
            begin
              reg654 <= reg656;
              reg655 = (($unsigned(forvar653[(3'h4):(3'h4)]) ?
                  wire646[(2'h2):(2'h2)] : $unsigned({(wire644 <<< reg654),
                      $unsigned(wire645)})) <= ((8'ha2) ^ reg651[(3'h5):(3'h4)]));
              reg659 = $signed((reg654 & $signed((~{(7'h44), (7'h43)}))));
            end
          if (reg659)
            begin
              reg660 = (~|((reg656[(3'h5):(1'h1)] ?
                      wire647[(3'h7):(3'h4)] : {$unsigned(wire645),
                          $signed((8'hb0))}) ?
                  wire649 : ($signed((&wire647)) ?
                      $signed(((8'hb9) ?
                          (7'h48) : reg656)) : ($signed(wire646) ?
                          (reg654 - reg653) : $unsigned(wire644)))));
              reg661 = wire652;
              reg662 = (((forvar653 ?
                      $unsigned($signed(wire647)) : ((reg654 ?
                              forvar653 : wire648) ?
                          $signed(forvar653) : forvar653[(2'h3):(1'h1)])) ^~ $signed(reg658)) ?
                  $unsigned((reg655 <= ({wire652, (8'hb7)} ~^ (reg660 ?
                      wire647 : reg653)))) : wire644[(1'h1):(1'h0)]);
              reg663 <= wire652;
              reg664 = $unsigned(reg659);
            end
          else
            begin
              reg660 = (|reg658);
              reg663 <= (^reg658);
              reg665 <= wire647[(3'h5):(1'h0)];
              reg666 <= reg663[(1'h0):(1'h0)];
            end
          if (wire646[(2'h3):(1'h0)])
            begin
              reg667 <= forvar653[(3'h4):(1'h1)];
              reg668 = $signed($unsigned($unsigned(($unsigned(wire646) ?
                  $signed(wire649) : (reg657 ^~ reg666)))));
              reg669 <= ($unsigned($signed((8'ha6))) >>> $signed($unsigned(((~|reg668) ?
                  (+(7'h46)) : (reg651 ? wire649 : reg662)))));
              reg670 <= (~^$unsigned((+reg651[(2'h2):(2'h2)])));
              reg671 = reg657;
            end
          else
            begin
              reg667 <= $unsigned(((reg658 || wire646) ?
                  $unsigned($signed((~^wire644))) : reg659[(5'h12):(5'h10)]));
            end
          for (forvar672 = (1'h0); (forvar672 < (3'h4)); forvar672 = (forvar672 + (1'h1)))
            begin
              reg673 = reg662[(4'hb):(3'h4)];
              reg674 = {($signed(($unsigned(reg656) ?
                      (reg654 >> wire646) : reg673[(4'hc):(4'ha)])) ^ {(~&{forvar672})})};
            end
          if ($unsigned({(+$unsigned(reg668))}))
            begin
              reg675 <= reg662[(4'he):(3'h6)];
              reg676 <= (-{($unsigned((reg657 ? reg666 : reg667)) - ({wire647,
                      reg661} <= {reg675}))});
              reg677 = wire645;
            end
          else
            begin
              reg677 = $unsigned((~^(!$unsigned((reg659 ? reg677 : reg659)))));
              reg678 <= (~^(-$unsigned({(reg674 ? reg676 : (8'ha8)),
                  (~&reg675)})));
              reg679 = $unsigned({reg654[(4'ha):(3'h4)]});
              reg680 = reg671[(3'h4):(2'h2)];
              reg681 <= (|$signed({{$unsigned(reg677)}}));
            end
        end
      if ($signed($unsigned((~^(^~(reg654 < reg667))))))
        begin
          reg682 <= (^~reg666[(4'he):(4'hc)]);
          for (forvar683 = (1'h0); (forvar683 < (2'h3)); forvar683 = (forvar683 + (1'h1)))
            begin
              reg684 = (7'h43);
            end
          for (forvar685 = (1'h0); (forvar685 < (3'h4)); forvar685 = (forvar685 + (1'h1)))
            begin
              reg686 <= (reg676 ?
                  $unsigned((~(^~reg674[(4'h8):(3'h7)]))) : $unsigned({$unsigned((reg674 ?
                          (8'haa) : forvar672))}));
              reg687 <= ($unsigned((reg679[(1'h1):(1'h0)] >> $unsigned(((7'h4a) ?
                      reg655 : reg676)))) ?
                  reg680 : reg677);
            end
          for (forvar688 = (1'h0); (forvar688 < (1'h1)); forvar688 = (forvar688 + (1'h1)))
            begin
              reg689 <= reg681;
              reg690 = $signed(({({reg660} != $signed(reg686))} <= (reg656 ?
                  ((reg665 <= reg678) ?
                      $signed(reg670) : $signed((8'h9d))) : (((8'hb7) ?
                      reg658 : wire646) < (wire644 >= reg662)))));
            end
        end
      else
        begin
          reg682 <= (wire646[(2'h2):(2'h2)] >= $signed(($signed($signed((8'hab))) > ((forvar653 ?
              wire646 : forvar653) << (!reg690)))));
          reg683 = $signed($unsigned((reg664 ?
              (reg654 ?
                  reg668[(5'h11):(5'h10)] : wire645[(2'h3):(1'h0)]) : (~^reg678))));
          reg684 = (&reg689[(3'h6):(3'h5)]);
          if (reg674)
            begin
              reg685 <= reg664[(3'h6):(3'h6)];
              reg688 = (~|forvar672[(3'h6):(1'h0)]);
              reg690 = $unsigned($unsigned({$signed((&reg680)),
                  ($signed(reg679) ?
                      forvar688[(2'h2):(2'h2)] : reg669[(3'h5):(1'h1)])}));
              reg691 <= {$unsigned(wire645), $signed(reg678)};
              reg692 = ({reg660[(1'h1):(1'h0)]} ?
                  reg673[(4'h9):(2'h2)] : {wire644});
            end
          else
            begin
              reg688 = reg686[(3'h5):(2'h2)];
              reg690 = (reg674[(4'hb):(1'h1)] >>> $unsigned((!{{reg651}})));
              reg692 = $signed((&$unsigned(reg667[(1'h1):(1'h1)])));
              reg693 <= $signed(($signed(reg653) ?
                  $signed($unsigned($signed(wire647))) : $signed((+(reg690 ?
                      reg662 : forvar683)))));
              reg694 = $signed((forvar653[(4'h8):(3'h6)] ?
                  wire648 : $signed(({reg675} == $unsigned((7'h42))))));
            end
          if ($signed(((&($unsigned((8'hba)) < $unsigned(reg691))) ?
              (7'h47) : reg690)))
            begin
              reg695 <= $unsigned(reg680);
              reg696 = reg682;
            end
          else
            begin
              reg696 = ((reg666[(4'hb):(1'h1)] ?
                      $unsigned($unsigned($unsigned(reg686))) : reg667[(3'h4):(2'h3)]) ?
                  (8'hb1) : ((((|reg665) ?
                          $unsigned(reg677) : $unsigned(reg657)) < $unsigned((reg666 <= reg664))) ?
                      {(wire649[(4'h9):(4'h9)] ?
                              forvar672[(2'h3):(1'h0)] : $signed((8'hb8)))} : (~(8'ha2))));
              reg697 = (8'hb0);
            end
        end
    end
  assign wire698 = $signed((reg651 ?
                       (^~(~^reg667[(1'h0):(1'h0)])) : {($signed(reg681) ^~ wire652[(4'ha):(3'h7)]),
                           ($signed(reg658) ?
                               (reg681 ? reg686 : reg681) : (~|reg675))}));
  assign wire699 = $unsigned((-(8'haa)));
  assign wire700 = (wire699 ^~ reg669[(2'h3):(2'h3)]);
  always
    @(posedge clk) begin
      if ((|(~(^~((reg667 ? (8'hb7) : reg686) ?
          (~reg657) : $unsigned(reg669))))))
        begin
          if ($signed(reg687[(1'h0):(1'h0)]))
            begin
              reg701 = $signed($unsigned((~^wire652)));
              reg702 = $unsigned((8'hb8));
              reg703 = $signed($unsigned($unsigned(($unsigned((8'ha8)) <= $unsigned(reg687)))));
              reg704 = reg686;
              reg705 = $signed((reg676 ?
                  (((reg691 ? reg695 : wire698) ?
                          reg665[(1'h0):(1'h0)] : $unsigned(reg702)) ?
                      (^~$signed((8'hbf))) : ({wire698, reg653} ?
                          wire648 : wire648[(3'h5):(3'h4)])) : $signed((wire646 ^ reg663))));
            end
          else
            begin
              reg701 = (((~|$unsigned(reg653)) < wire652) > (!(^~$signed(reg665[(4'hb):(3'h6)]))));
              reg706 <= reg653;
              reg707 = reg667[(3'h4):(1'h0)];
            end
          reg708 = (7'h42);
          reg709 <= (reg704[(3'h4):(3'h4)] || {wire646});
          if (reg658)
            begin
              reg710 <= reg701;
              reg711 = $unsigned(($unsigned(reg653) - (|($signed(wire648) + (reg651 ?
                  reg678 : reg658)))));
              reg712 <= $signed($unsigned($unsigned(reg703)));
              reg713 = (&$signed({(~|(reg667 ? reg708 : reg657)),
                  (reg707 * reg658)}));
            end
          else
            begin
              reg710 <= $unsigned(reg653);
              reg711 = ((((reg670[(3'h6):(3'h6)] ?
                          wire699 : {reg676,
                              (8'hb4)}) - (reg712[(3'h7):(1'h0)] << reg713[(4'ha):(3'h4)])) ?
                      $signed($signed($unsigned(reg705))) : (((reg703 && reg709) <<< (~^reg667)) - (!(8'h9c)))) ?
                  (!(((reg654 <= reg657) ?
                      (8'hb8) : wire699) & reg687)) : ((8'ha7) ?
                      {((&reg695) && $signed(reg695)),
                          (((7'h44) >= reg709) ?
                              reg687 : $unsigned(wire648))} : $signed((reg713 ?
                          (reg691 ? wire646 : reg712) : {reg685}))));
              reg712 <= ((-reg685) ?
                  (-reg712) : ($signed(reg658[(1'h0):(1'h0)]) | $unsigned((wire652[(5'h12):(4'hd)] >>> (|wire698)))));
              reg713 = ({reg701[(4'he):(4'h9)]} ?
                  ($unsigned($unsigned((+wire652))) ?
                      (($signed(reg711) ?
                              (reg709 && (8'h9e)) : $unsigned(reg708)) ?
                          reg657 : {$signed(reg653),
                              (~^(8'ha5))}) : ((-{reg702}) <= $signed(reg691[(3'h5):(3'h4)]))) : ((reg701 + (|$unsigned(reg676))) || wire644));
            end
          reg714 <= ((8'hab) < (8'hae));
        end
      else
        begin
          reg706 <= $unsigned(reg685[(4'hb):(4'h9)]);
          reg707 = reg687;
          reg709 <= $unsigned({$signed(reg676[(3'h4):(2'h3)])});
        end
      reg715 <= ($unsigned(wire699) == $unsigned((((wire645 ~^ reg710) ?
              {reg663, reg667} : (~&reg705)) ?
          {reg685, (|reg665)} : ((reg713 != reg709) <<< (reg657 ?
              reg701 : reg712)))));
      if ($unsigned(((^~(7'h44)) >= {$signed($unsigned(reg669)),
          (+reg657[(3'h5):(2'h2)])})))
        begin
          reg716 <= (8'hba);
          for (forvar717 = (1'h0); (forvar717 < (3'h4)); forvar717 = (forvar717 + (1'h1)))
            begin
              reg718 <= $signed(reg715[(3'h7):(1'h0)]);
            end
          for (forvar719 = (1'h0); (forvar719 < (2'h3)); forvar719 = (forvar719 + (1'h1)))
            begin
              reg720 <= ((|$unsigned((reg675[(3'h7):(2'h3)] & ((8'hb1) && reg682)))) ?
                  ($unsigned(reg686) != ({wire699[(2'h3):(2'h3)],
                      $signed(reg702)} ^ reg657[(3'h5):(1'h0)])) : ($signed(($signed(reg686) ?
                      $signed(reg707) : ((8'hb3) ?
                          reg715 : reg702))) >> {({(7'h41),
                          wire700} ~^ {reg665})}));
              reg721 = (reg706[(4'h9):(4'h8)] ?
                  $unsigned($signed((!(reg670 ?
                      reg711 : reg705)))) : (-reg701[(4'hf):(4'h9)]));
              reg722 <= $unsigned(reg676[(1'h1):(1'h0)]);
              reg723 <= {((~($unsigned(wire700) ?
                      $signed(reg666) : {reg676})) >> reg706),
                  (reg676[(1'h1):(1'h0)] ?
                      {(!(reg675 ? reg708 : wire645)),
                          (^(~&wire647))} : $unsigned((^wire699[(4'h8):(4'h8)])))};
            end
        end
      else
        begin
          reg717 = reg658;
          for (forvar718 = (1'h0); (forvar718 < (2'h2)); forvar718 = (forvar718 + (1'h1)))
            begin
              reg719 <= {$unsigned(reg701)};
            end
          for (forvar720 = (1'h0); (forvar720 < (2'h2)); forvar720 = (forvar720 + (1'h1)))
            begin
              reg721 = (($signed($unsigned((reg721 ? reg669 : forvar719))) ?
                  ((~&$unsigned(reg723)) ?
                      reg719 : ($signed((8'h9e)) * $unsigned((8'ha7)))) : (reg686 ?
                      {$signed(reg704), (^(8'h9d))} : (~&reg689))) >= wire699);
              reg722 <= $signed((|$unsigned(((^~reg675) ?
                  (wire647 <= (7'h4a)) : (reg716 ? reg701 : reg721)))));
              reg723 <= ($unsigned(reg676) != (reg656[(3'h5):(1'h1)] ?
                  reg723[(4'hb):(1'h0)] : reg706[(1'h0):(1'h0)]));
            end
          reg724 = ((~$signed((reg714[(3'h7):(3'h5)] ?
              (!reg665) : ((8'ha7) + reg686)))) && (reg691[(1'h0):(1'h0)] * $signed((reg723[(4'he):(4'hb)] ?
              (reg669 == reg704) : wire699))));
          if ((((~$unsigned((wire645 - wire698))) ?
                  $unsigned($signed((reg703 + reg720))) : forvar719[(1'h1):(1'h0)]) ?
              ($unsigned(forvar717[(3'h4):(1'h1)]) ?
                  {$unsigned((~reg669))} : $signed(wire647)) : (~^$signed(reg691[(2'h3):(1'h0)]))))
            begin
              reg725 <= $signed((($signed((reg678 ?
                      reg669 : reg681)) & {(+wire647)}) ?
                  reg654[(1'h1):(1'h1)] : (!reg702[(1'h0):(1'h0)])));
              reg726 <= $signed((($signed(wire648) == wire652) ?
                  (8'h9d) : $unsigned(((!reg724) ?
                      $signed(reg681) : (-reg719)))));
              reg727 = $unsigned(reg717[(3'h7):(2'h2)]);
              reg728 <= reg667[(1'h0):(1'h0)];
              reg729 = ({forvar717,
                  (reg654 ?
                      $unsigned(reg670) : (-reg714))} > {((-((8'hbd) || reg669)) ?
                      (~&(~&reg721)) : $signed({reg727, reg651})),
                  $unsigned(((^~forvar720) || (reg682 >= wire646)))});
            end
          else
            begin
              reg727 = reg725;
              reg728 <= ((reg725[(1'h1):(1'h0)] ?
                      $unsigned({$unsigned((7'h49))}) : (reg682 ~^ $signed((reg705 ?
                          reg665 : reg714)))) ?
                  $signed((($signed(reg719) ^ (reg691 ? reg716 : wire699)) ?
                      $signed($signed(forvar718)) : ($unsigned(forvar720) == {(8'hb3),
                          reg729}))) : (($unsigned(reg709[(4'hd):(3'h6)]) << $unsigned(reg695)) << (!$signed($signed(wire649)))));
            end
        end
      for (forvar730 = (1'h0); (forvar730 < (1'h0)); forvar730 = (forvar730 + (1'h1)))
        begin
          for (forvar731 = (1'h0); (forvar731 < (1'h1)); forvar731 = (forvar731 + (1'h1)))
            begin
              reg732 = wire700[(4'h9):(2'h3)];
            end
        end
      if ($unsigned(($signed(reg665[(1'h0):(1'h0)]) ?
          reg670[(4'hf):(4'h8)] : reg669)))
        begin
          for (forvar733 = (1'h0); (forvar733 < (3'h4)); forvar733 = (forvar733 + (1'h1)))
            begin
              reg734 = reg667[(2'h2):(1'h0)];
              reg735 = ({(~&$unsigned({reg707}))} ?
                  ($signed((^reg681[(3'h4):(1'h1)])) ?
                      reg651 : (wire645 ? reg725 : wire700)) : reg720);
            end
          for (forvar736 = (1'h0); (forvar736 < (2'h2)); forvar736 = (forvar736 + (1'h1)))
            begin
              reg737 <= (~&($signed((~&$unsigned(reg687))) ?
                  (((reg667 ?
                      reg711 : forvar717) ~^ reg711[(2'h3):(2'h2)]) >>> ((reg710 * forvar736) << wire647[(3'h7):(2'h3)])) : (~^reg666)));
              reg738 <= (^(^~reg656[(4'h8):(1'h1)]));
              reg739 = reg653;
              reg740 = $unsigned((|reg715[(3'h4):(1'h1)]));
            end
        end
      else
        begin
          reg733 = (reg712 ? $signed((!reg724)) : $unsigned(reg670));
          reg736 <= reg713;
          if ((($unsigned($unsigned(reg653[(3'h5):(1'h0)])) > ($unsigned($signed(reg669)) ?
                  $signed($signed(reg739)) : {$signed((7'h44))})) ?
              reg656[(3'h6):(2'h2)] : reg705))
            begin
              reg737 <= (((~&$unsigned(((7'h49) ? reg657 : reg709))) ?
                      (+(~|(reg682 - (7'h49)))) : (8'hbf)) ?
                  ((reg734[(1'h1):(1'h0)] ?
                      (&reg693) : reg665[(4'h9):(3'h7)]) >> reg705) : (!(!(reg714[(2'h2):(1'h0)] + (-wire644)))));
              reg738 <= ((($unsigned($unsigned(reg663)) ?
                      reg656[(2'h2):(2'h2)] : $signed(reg702[(4'ha):(4'ha)])) ?
                  (&(reg738 >>> {reg657,
                      (8'had)})) : $signed(reg717)) - {($signed($signed(reg725)) ?
                      $unsigned((|(8'ha9))) : (^~wire652[(4'h8):(2'h3)])),
                  $signed((&(reg719 ? reg722 : (8'hb5))))});
              reg741 <= reg666[(3'h6):(2'h3)];
              reg742 = (|(|reg658[(1'h1):(1'h1)]));
              reg743 <= reg721[(4'h9):(1'h1)];
            end
          else
            begin
              reg739 = ((((wire645 <<< (^~reg653)) + {reg726}) ?
                      ((reg712[(4'hd):(3'h5)] >> {reg695, wire648}) ?
                          (~^$signed(reg733)) : reg707[(3'h4):(2'h2)]) : (reg721 & ((reg708 ?
                          reg691 : (8'haf)) > (reg657 >>> reg676)))) ?
                  reg667 : reg657);
              reg741 <= {forvar731[(3'h5):(3'h5)],
                  ((($signed(reg702) ~^ (reg670 ?
                      reg736 : (8'h9d))) >> ((&reg708) != (^~reg705))) <<< (reg726 ^~ reg720))};
              reg742 = $signed($signed(reg738[(1'h0):(1'h0)]));
              reg743 <= $signed(((!$signed($unsigned(wire647))) * reg676));
              reg744 = reg707;
            end
          for (forvar745 = (1'h0); (forvar745 < (2'h2)); forvar745 = (forvar745 + (1'h1)))
            begin
              reg746 = (!(reg709 ? reg734 : $signed((reg717 ^ reg737))));
              reg747 = reg678[(3'h7):(3'h5)];
            end
        end
    end
  always
    @(posedge clk) begin
      if ((~|$signed(reg719)))
        begin
          reg748 = $signed(wire645[(4'h8):(3'h4)]);
          for (forvar749 = (1'h0); (forvar749 < (2'h2)); forvar749 = (forvar749 + (1'h1)))
            begin
              reg750 = reg678;
              reg751 = {{($signed((~^reg743)) ?
                          reg669[(3'h5):(1'h0)] : {wire645[(2'h2):(1'h0)],
                              (reg706 >= (8'hab))})},
                  $signed(($unsigned($signed(reg658)) ? reg669 : reg720))};
              reg752 <= (~&$signed(({(|wire648)} ?
                  (^(8'ha0)) : (reg665 ~^ $unsigned(reg723)))));
              reg753 <= $signed(((-reg693) >= $unsigned(((reg686 ?
                      reg689 : reg709) ?
                  $unsigned((8'hb2)) : $unsigned(reg719)))));
              reg754 <= {$signed((wire648[(3'h6):(1'h1)] ?
                      (~^$signed(reg658)) : (!$unsigned(reg753))))};
            end
        end
      else
        begin
          for (forvar748 = (1'h0); (forvar748 < (1'h1)); forvar748 = (forvar748 + (1'h1)))
            begin
              reg749 = ($signed(reg725[(2'h3):(2'h2)]) | $signed($unsigned((reg663 >>> $unsigned(reg720)))));
              reg752 <= $signed(reg685);
              reg753 <= $unsigned(($signed(reg666) ?
                  $signed(({(7'h46)} ?
                      reg658[(3'h6):(2'h3)] : reg754[(5'h13):(3'h5)])) : ({reg706[(1'h0):(1'h0)]} != ((+wire647) < (reg710 ?
                      reg695 : reg715)))));
              reg754 <= (^$signed((reg653 != $signed(reg715))));
              reg755 <= (({(!{reg685, reg687})} || (((wire644 ?
                  (8'hb3) : reg752) - $unsigned(reg687)) < (reg715[(4'h9):(4'h9)] ?
                  ((8'ha0) >> reg728) : $signed(wire644)))) < $signed((reg667 != reg676[(3'h7):(3'h4)])));
            end
        end
      if ($signed({($signed(reg743[(4'he):(4'hd)]) ?
              (&reg689[(1'h0):(1'h0)]) : reg693[(1'h1):(1'h1)])}))
        begin
          reg756 = reg653[(3'h7):(3'h5)];
          reg757 <= $unsigned(((($unsigned(reg689) >>> (7'h48)) ?
              ($signed(reg687) ?
                  reg675[(2'h2):(1'h1)] : $signed(reg725)) : (&(~^reg716))) > $signed(reg750[(1'h1):(1'h1)])));
          reg758 <= (reg714[(1'h1):(1'h0)] ?
              reg695[(1'h0):(1'h0)] : $signed(reg751[(2'h2):(2'h2)]));
        end
      else
        begin
          reg756 = $signed(reg657[(3'h6):(1'h0)]);
          for (forvar757 = (1'h0); (forvar757 < (2'h2)); forvar757 = (forvar757 + (1'h1)))
            begin
              reg759 = {$unsigned(reg756[(4'ha):(1'h0)]),
                  {$unsigned((+(7'h42)))}};
              reg760 <= reg710;
              reg761 <= ($unsigned((reg725[(3'h5):(3'h4)] != (~^$unsigned(reg718)))) ?
                  reg657 : (-reg756[(3'h4):(2'h2)]));
              reg762 <= (~|reg754);
            end
          reg763 = $signed((($signed((reg712 != reg728)) || reg682[(1'h0):(1'h0)]) ?
              {$unsigned($unsigned(reg749)),
                  ($unsigned(reg715) ?
                      (~&reg718) : (reg706 + reg665))} : (reg723[(3'h4):(2'h2)] >= $unsigned((~reg741)))));
          for (forvar764 = (1'h0); (forvar764 < (2'h3)); forvar764 = (forvar764 + (1'h1)))
            begin
              reg765 <= (~|($unsigned(((+(8'ha2)) ?
                  reg681[(5'h11):(3'h7)] : (-reg686))) ^ (^~reg743)));
              reg766 = ({$signed($unsigned((~&reg712))),
                  ((^~$unsigned(reg763)) ?
                      {$unsigned(reg765),
                          $signed(reg675)} : $signed(wire646[(2'h2):(1'h0)]))} && {reg710[(2'h2):(1'h1)],
                  wire699});
              reg767 <= wire699;
              reg768 <= (((^~($signed((8'hb5)) + (reg682 ?
                      (8'hbf) : (8'hb7)))) <= reg765) ?
                  ($signed($signed((~^reg709))) ?
                      ($unsigned(reg686) ^~ $signed($unsigned((8'hb3)))) : reg689[(1'h0):(1'h0)]) : (|(({reg748} ?
                          reg743 : $signed(reg765)) ?
                      $signed($signed(reg654)) : reg720)));
              reg769 <= $signed((~(|{(^reg709)})));
            end
        end
    end
  always
    @(posedge clk) begin
      for (forvar770 = (1'h0); (forvar770 < (2'h3)); forvar770 = (forvar770 + (1'h1)))
        begin
          reg771 = ($unsigned((reg691 | $signed((reg654 ? reg665 : reg658)))) ?
              ({(reg720[(1'h0):(1'h0)] <= $unsigned(wire698)),
                  ((reg726 | reg678) ?
                      (&reg663) : reg657[(1'h0):(1'h0)])} ~^ $signed(reg651)) : $unsigned($signed((-(reg676 ?
                  reg765 : (8'ha6))))));
          if (((~($signed($signed(wire647)) | (reg765[(4'h9):(1'h1)] - $signed(reg693)))) ?
              reg651 : (~reg670)))
            begin
              reg772 <= reg723;
            end
          else
            begin
              reg772 <= ($signed($signed($unsigned(reg651))) - reg736);
              reg773 = ((~&reg670[(3'h6):(3'h4)]) != ($signed(reg771) ?
                  reg715 : ((|$signed(reg728)) << $unsigned((8'haa)))));
              reg774 = ($signed(wire700[(2'h3):(1'h0)]) ^~ reg772[(1'h0):(1'h0)]);
              reg775 = (($signed($signed(wire698[(4'h8):(2'h2)])) && $signed(((~&reg755) ?
                      {reg722} : reg752))) ?
                  $signed(((^reg710[(2'h2):(1'h1)]) ?
                      $signed({reg754}) : $unsigned(wire648[(5'h11):(2'h3)]))) : (reg657 & $unsigned(((reg675 ?
                          wire699 : wire644) ?
                      {reg773} : $signed(reg762)))));
            end
          for (forvar776 = (1'h0); (forvar776 < (2'h3)); forvar776 = (forvar776 + (1'h1)))
            begin
              reg777 <= ($unsigned((~&((~&reg651) <<< $unsigned(reg670)))) ?
                  (~reg718[(5'h14):(1'h1)]) : (~(($unsigned(reg738) >> reg712[(4'h8):(3'h6)]) ?
                      $signed((8'hb7)) : (reg723 > (reg657 != wire646)))));
              reg778 = (((reg743[(4'hc):(4'h9)] ?
                      wire645 : (!(reg685 ? reg737 : (8'hb5)))) ?
                  $signed(reg695) : ($signed((reg719 ^~ (7'h45))) && ($unsigned(wire649) * {reg761}))) >> {(reg773[(4'h9):(4'h8)] >= ((reg755 ?
                          (8'hb8) : reg687) ?
                      $unsigned(reg709) : $unsigned(wire652)))});
              reg779 <= (-(~&reg686));
              reg780 = (!reg718);
              reg781 = (-((reg718[(5'h15):(4'hc)] <<< (+(|(8'ha9)))) >>> $signed(reg736)));
            end
          for (forvar782 = (1'h0); (forvar782 < (1'h1)); forvar782 = (forvar782 + (1'h1)))
            begin
              reg783 = reg657[(2'h2):(2'h2)];
              reg784 <= (((~reg695) != reg783) || $unsigned({(^~(reg736 || reg656))}));
            end
        end
      if (reg725[(1'h0):(1'h0)])
        begin
          for (forvar785 = (1'h0); (forvar785 < (1'h1)); forvar785 = (forvar785 + (1'h1)))
            begin
              reg786 <= reg762[(3'h5):(1'h0)];
              reg787 = {reg775};
              reg788 <= $signed(($unsigned((^(|reg669))) | $unsigned((~|reg778))));
              reg789 <= reg787;
            end
          if ((($unsigned(reg710) ?
                  {((reg657 ? reg758 : reg761) ?
                          reg761[(4'he):(4'hb)] : $signed((8'hab)))} : ($unsigned($unsigned(reg779)) ?
                      (reg693 >= $signed(wire700)) : $unsigned((reg774 == reg719)))) ?
              $signed($signed($unsigned($signed(reg651)))) : $signed((~|(-(~&reg755))))))
            begin
              reg790 <= reg736;
              reg791 <= (8'hbf);
              reg792 <= (reg666[(1'h0):(1'h0)] ?
                  $signed((~|$signed(reg712))) : ({reg653} != {$signed((^wire646)),
                      $signed((&(8'ha2)))}));
            end
          else
            begin
              reg793 = ((reg777 == ($unsigned((8'ha4)) ?
                  ((+wire646) | $signed(forvar770)) : {wire647,
                      (reg752 ?
                          reg691 : wire648)})) ~^ (!reg768[(3'h6):(1'h0)]));
              reg794 <= $unsigned(((!reg691[(4'h8):(3'h5)]) | (reg710[(1'h1):(1'h1)] ?
                  ($signed(reg780) ^ (reg738 < reg695)) : {$unsigned(reg765),
                      wire644})));
            end
        end
      else
        begin
          if ({$unsigned(($unsigned(wire700) ?
                  wire646[(2'h2):(1'h0)] : ((reg687 ? reg709 : reg783) ?
                      (reg762 - (8'h9e)) : $signed((8'hb8))))),
              $unsigned(wire652[(4'h9):(3'h7)])})
            begin
              reg785 <= {($unsigned(({reg712} ?
                          reg669 : reg793[(4'h9):(1'h1)])) ?
                      (|(^(^(8'hb0)))) : ((~^(reg761 ? reg768 : forvar776)) ?
                          reg757 : forvar776)),
                  (&reg755)};
              reg786 <= (^~{$signed(reg669)});
              reg788 <= $unsigned($unsigned((7'h4a)));
              reg793 = reg653;
              reg795 = (~reg743[(3'h6):(3'h6)]);
            end
          else
            begin
              reg785 <= (reg777[(2'h2):(2'h2)] ?
                  reg752[(1'h0):(1'h0)] : $unsigned({(+(^(7'h46)))}));
              reg786 <= (^$unsigned(reg669[(1'h1):(1'h0)]));
              reg787 = (~$signed($signed((reg761[(3'h7):(1'h1)] ?
                  (!wire700) : (reg738 ? reg788 : forvar770)))));
              reg793 = ($unsigned((~&$unsigned(reg720))) < reg714[(4'hb):(4'h8)]);
            end
          for (forvar796 = (1'h0); (forvar796 < (1'h1)); forvar796 = (forvar796 + (1'h1)))
            begin
              reg797 = reg691;
              reg798 = ((reg787[(1'h1):(1'h1)] ?
                      $signed(({reg783} > $signed(reg676))) : {$signed($signed(reg778)),
                          ($signed(reg757) ?
                              (^~reg778) : (forvar782 ? wire647 : wire645))}) ?
                  ((((reg714 ~^ reg793) << $signed(reg682)) >> reg691) ?
                      (^~(~(reg706 >>> reg774))) : $unsigned(forvar782)) : $signed($unsigned(($signed(reg792) ^ $unsigned((7'h48))))));
              reg799 = (~^(~|(7'h46)));
              reg800 <= ($unsigned(reg790[(2'h2):(1'h0)]) < (reg761 ~^ $unsigned(reg726[(4'hb):(4'h8)])));
            end
          if (reg653)
            begin
              reg801 = $signed(((8'hb0) ?
                  ($unsigned({(8'haa),
                      reg710}) > (^~$signed(forvar782))) : (($signed(reg716) ?
                      {reg777, (8'ha4)} : $unsigned(reg737)) || reg762)));
              reg802 = ((($signed((~&reg791)) < (~^(reg773 ?
                          reg687 : wire699))) ?
                      ((~^$unsigned(reg794)) ?
                          (7'h48) : $signed({reg800, reg689})) : ((reg666 ?
                          $signed(reg771) : (reg777 ?
                              reg656 : wire645)) == {reg738, reg653})) ?
                  {(+((reg801 && wire698) & (reg710 ^ reg736))),
                      {reg784[(1'h1):(1'h0)],
                          {reg795}}} : $unsigned({$unsigned(reg654[(3'h4):(1'h0)])}));
            end
          else
            begin
              reg803 <= $signed((reg725[(1'h1):(1'h0)] != reg758));
              reg804 <= (wire648 ? $unsigned(reg795[(4'hf):(3'h7)]) : reg736);
            end
          reg805 <= reg788[(4'hc):(3'h7)];
        end
      reg806 <= reg676;
      reg807 <= reg758;
      for (forvar808 = (1'h0); (forvar808 < (2'h3)); forvar808 = (forvar808 + (1'h1)))
        begin
          for (forvar809 = (1'h0); (forvar809 < (1'h1)); forvar809 = (forvar809 + (1'h1)))
            begin
              reg810 <= $signed((~&wire649));
              reg811 = reg753;
            end
          reg812 <= ({$signed((7'h46))} < (($unsigned($unsigned(reg695)) ?
              ($signed((8'hb7)) && $unsigned(forvar782)) : (&$signed(reg725))) ^ (~&reg760[(2'h3):(2'h2)])));
          if (reg654)
            begin
              reg813 <= ($unsigned(reg755) ?
                  ((&{reg798}) ?
                      (reg691 ?
                          wire644 : ((reg743 ?
                              reg681 : forvar782) >= reg693[(2'h3):(1'h0)])) : $signed({reg710})) : $unsigned(reg804[(4'hd):(2'h3)]));
              reg814 <= $unsigned($unsigned($signed(reg687)));
              reg815 <= {((~((reg725 << reg806) ? reg737 : $signed(wire645))) ?
                      $signed($signed(((8'hb8) ? reg779 : (7'h46)))) : (reg788 ?
                          (~&{(8'h9c)}) : reg797[(4'h9):(4'h9)]))};
              reg816 = {($unsigned($unsigned($unsigned(reg791))) >> reg807),
                  reg773};
            end
          else
            begin
              reg813 <= (-(~&(((&reg720) ?
                  (wire644 == reg780) : reg755[(1'h0):(1'h0)]) << ($unsigned((8'hb8)) ?
                  ((8'h9e) | (8'hbd)) : (reg755 ? (8'hb4) : reg710)))));
              reg816 = $unsigned((~reg675));
            end
          reg817 <= {$unsigned($signed(reg761[(1'h1):(1'h0)])),
              ({reg728} ^ $signed($unsigned($unsigned(reg780))))};
          reg818 = reg786;
        end
    end
  always
    @(posedge clk) begin
      if ($unsigned(((reg815[(3'h6):(3'h5)] >> (8'hb6)) << $unsigned(reg728[(2'h3):(1'h1)]))))
        begin
          reg819 = (($unsigned(((~|reg803) || {reg665})) ?
              $unsigned(($signed(reg719) * reg769[(5'h10):(1'h0)])) : (~|(reg709 < {reg772}))) < (($unsigned((+reg658)) == $unsigned((reg656 | reg686))) <<< (~^({reg653,
                  reg758} ?
              (reg685 <<< reg725) : reg726[(4'h8):(3'h6)]))));
          for (forvar820 = (1'h0); (forvar820 < (1'h1)); forvar820 = (forvar820 + (1'h1)))
            begin
              reg821 <= (^~{(reg720[(2'h2):(1'h1)] ?
                      $signed(reg719) : (wire652 & $signed(reg725))),
                  ((~^reg817) * (~&(reg736 && reg738)))});
              reg822 <= (~^reg767);
              reg823 = reg814[(5'h11):(4'ha)];
            end
          reg824 <= $unsigned(reg772[(2'h3):(2'h3)]);
          for (forvar825 = (1'h0); (forvar825 < (1'h0)); forvar825 = (forvar825 + (1'h1)))
            begin
              reg826 = $signed($signed((reg736 <<< (^$signed(reg685)))));
              reg827 = (($unsigned(reg794[(5'h14):(2'h2)]) ?
                      $signed($unsigned((^~reg667))) : $signed($unsigned($signed(reg779)))) ?
                  (|$signed((~&reg710))) : $unsigned(reg762));
              reg828 <= reg669;
              reg829 <= $unsigned((8'hb8));
              reg830 <= ((^$unsigned(reg760[(3'h5):(1'h0)])) == ((reg693 ?
                      ($signed(reg687) ?
                          {(8'hac)} : reg803) : $signed($unsigned(reg760))) ?
                  (reg817[(4'hd):(3'h7)] ?
                      reg736[(1'h0):(1'h0)] : (7'h41)) : ((&$unsigned(reg726)) ?
                      wire698[(3'h4):(2'h2)] : forvar825[(3'h6):(3'h5)])));
            end
          for (forvar831 = (1'h0); (forvar831 < (2'h2)); forvar831 = (forvar831 + (1'h1)))
            begin
              reg832 <= $signed(reg791[(3'h5):(1'h1)]);
              reg833 <= reg738;
              reg834 = (reg805[(3'h5):(1'h1)] ?
                  $signed((wire648 ?
                      ((-reg678) ?
                          (|reg710) : {reg813}) : forvar820)) : (~&reg789[(3'h5):(2'h3)]));
              reg835 = ((!reg790[(4'hb):(3'h7)]) ?
                  ((+(reg712 || $unsigned(wire700))) == $signed((reg779 + $signed(reg738)))) : reg830);
              reg836 <= $signed(reg784[(3'h4):(3'h4)]);
            end
        end
      else
        begin
          reg819 = reg804[(4'hf):(4'hc)];
          reg820 <= ((8'ha6) && $unsigned((8'hab)));
          for (forvar821 = (1'h0); (forvar821 < (1'h0)); forvar821 = (forvar821 + (1'h1)))
            begin
              reg822 <= reg800[(2'h2):(1'h1)];
              reg823 = {{$unsigned({(forvar820 ? (8'h9e) : reg669)})},
                  ($unsigned(($unsigned(reg743) ^~ ((8'ha9) != (8'ha8)))) ?
                      ((+$signed(reg755)) ?
                          $unsigned((reg758 ?
                              reg785 : (8'hb5))) : $unsigned(wire649)) : (^reg753))};
              reg825 = (8'ha6);
              reg828 <= ((8'hb0) & $unsigned($unsigned(($unsigned(reg653) ?
                  reg685 : reg682[(2'h2):(1'h1)]))));
            end
        end
      for (forvar837 = (1'h0); (forvar837 < (2'h3)); forvar837 = (forvar837 + (1'h1)))
        begin
          for (forvar838 = (1'h0); (forvar838 < (2'h2)); forvar838 = (forvar838 + (1'h1)))
            begin
              reg839 <= (((!wire646[(2'h2):(1'h0)]) ? reg833 : reg657) ?
                  reg718[(4'hc):(4'h8)] : $unsigned(reg830));
              reg840 = (!($signed(wire652[(5'h14):(5'h11)]) ?
                  reg657[(3'h5):(3'h4)] : {$signed(reg827[(1'h0):(1'h0)])}));
              reg841 <= ($signed(reg828[(2'h2):(1'h0)]) | ($unsigned($signed({reg670})) - reg814));
            end
          reg842 = $unsigned(reg758[(5'h12):(3'h7)]);
          reg843 = $unsigned((~|$unsigned($unsigned($unsigned(reg836)))));
        end
    end
  assign wire844 = $signed($unsigned(((-{(8'ha8), reg658}) ?
                       ((-reg718) & reg829) : $unsigned((~&(8'h9c))))));
  assign wire845 = reg772[(2'h3):(1'h1)];
  always
    @(posedge clk) begin
      if (reg757[(2'h3):(1'h1)])
        begin
          reg846 = reg753[(3'h4):(2'h2)];
          reg847 <= reg839[(2'h2):(1'h0)];
          for (forvar848 = (1'h0); (forvar848 < (1'h0)); forvar848 = (forvar848 + (1'h1)))
            begin
              reg849 <= (((({reg715} ?
                      {reg682,
                          reg791} : $unsigned(wire845)) > ({reg810} >= (reg719 ?
                      reg807 : reg653))) ?
                  reg804[(3'h5):(3'h4)] : ({reg653[(1'h0):(1'h0)],
                          (reg769 ? (7'h44) : reg765)} ?
                      (((8'hb9) || reg800) & wire844[(5'h16):(4'hb)]) : $signed($unsigned(reg738)))) <= ((reg777[(4'h8):(2'h3)] ^ $unsigned({wire652})) ?
                  (^{$signed(reg753),
                      reg719[(2'h3):(2'h3)]}) : (&({reg803} ^ $signed(reg803)))));
            end
          if (reg691)
            begin
              reg850 = {($unsigned(($signed(reg803) ?
                      reg821 : (|(8'ha1)))) || (!$unsigned(reg715[(3'h7):(3'h5)])))};
              reg851 = $unsigned((reg695[(1'h1):(1'h0)] ?
                  reg841[(3'h6):(2'h3)] : {reg788,
                      (reg719[(2'h3):(1'h0)] - reg830)}));
              reg852 = (8'hb3);
              reg853 <= wire652;
              reg854 <= ({(8'hbd)} ?
                  $signed(reg714[(3'h5):(1'h1)]) : (($signed($signed(reg682)) ?
                          (reg669 ?
                              wire647 : (wire644 ^~ reg654)) : reg846[(3'h4):(1'h1)]) ?
                      reg788[(3'h5):(2'h2)] : (($unsigned(reg653) ?
                          (8'hb7) : $unsigned((8'ha1))) == (reg792[(1'h0):(1'h0)] <= reg665))));
            end
          else
            begin
              reg853 <= ($signed((~^{$unsigned(reg761)})) ?
                  reg681[(3'h5):(3'h4)] : $unsigned(reg805));
              reg855 = (reg722[(3'h6):(3'h5)] | reg687);
              reg856 <= reg728[(1'h1):(1'h1)];
              reg857 <= {((wire649[(3'h6):(1'h1)] > {(reg758 && reg726),
                          (reg761 ? wire700 : reg653)}) ?
                      (&(-{reg786})) : (($unsigned(reg815) >> (|reg836)) ?
                          (&reg847) : ({reg709, reg754} ?
                              (~reg754) : (reg761 << reg725))))};
            end
          reg858 = $unsigned((|(&(~|(reg665 * reg836)))));
        end
      else
        begin
          if ((($signed($signed((reg849 ?
                  (8'hae) : reg737))) - $signed(reg726[(3'h5):(3'h5)])) ?
              reg858 : $unsigned(reg681)))
            begin
              reg846 = (((~|((reg768 ? reg854 : reg761) ?
                      {reg691, reg856} : (~&reg682))) ?
                  $unsigned(((!wire699) ?
                      (&(8'hb0)) : {reg678,
                          wire699})) : $signed(reg718)) & $signed(reg841[(5'h14):(4'ha)]));
              reg848 = $signed({reg725[(3'h4):(2'h3)], reg757[(4'hb):(2'h2)]});
              reg849 <= ((reg829 == $unsigned(reg760[(1'h0):(1'h0)])) ?
                  $signed((!((!reg695) ?
                      reg857 : (reg736 ^ reg794)))) : $signed({((reg657 && reg667) >> $unsigned(wire700))}));
            end
          else
            begin
              reg847 <= ($signed({reg675[(3'h5):(1'h1)]}) != ($signed(reg741[(2'h2):(1'h1)]) ?
                  reg839[(3'h4):(1'h0)] : (^~(8'hb8))));
              reg849 <= (reg712 ? $unsigned(reg792) : wire649);
            end
          reg850 = reg689;
          reg851 = (^{$signed((((8'hbe) ?
                  (7'h47) : reg754) <<< reg784[(3'h5):(1'h1)])),
              (^({reg738} << (reg682 > (8'haa))))});
          reg852 = $unsigned(($signed({reg815[(4'ha):(4'h9)],
              $signed(reg681)}) ~^ (~|$signed((wire699 && reg850)))));
        end
      reg859 = (7'h41);
      for (forvar860 = (1'h0); (forvar860 < (2'h2)); forvar860 = (forvar860 + (1'h1)))
        begin
          reg861 = reg804;
          for (forvar862 = (1'h0); (forvar862 < (2'h3)); forvar862 = (forvar862 + (1'h1)))
            begin
              reg863 = $signed($signed($signed((^~$unsigned(reg804)))));
              reg864 = reg678;
              reg865 = (!{$signed(($unsigned(reg669) | {reg710})),
                  $signed((reg676[(1'h1):(1'h0)] - ((8'hac) >> (7'h43))))});
              reg866 <= reg685[(4'he):(3'h7)];
              reg867 = reg794;
            end
        end
      reg868 = reg752;
      reg869 <= reg786;
    end
  assign wire870 = $unsigned($signed($unsigned((!reg752))));
  always
    @(posedge clk) begin
      reg871 <= $unsigned((($signed(reg686) ?
          ((!reg822) >= $unsigned((8'h9c))) : {reg836}) ^~ (reg714[(3'h6):(3'h4)] ?
          ((reg738 ? reg685 : reg830) & (|reg657)) : $unsigned((^reg741)))));
      reg872 = (wire652[(2'h2):(2'h2)] & reg723[(4'hc):(1'h1)]);
    end
  always
    @(posedge clk) begin
      if ({reg790})
        begin
          reg873 <= reg658;
          if (((reg789[(3'h5):(1'h0)] ?
              ($unsigned($unsigned(reg777)) ?
                  ((reg854 & reg653) ^ $unsigned(reg856)) : reg686[(2'h3):(2'h3)]) : reg693) ^ ((-reg806[(3'h4):(1'h1)]) ?
              $signed($unsigned(reg792)) : $unsigned({(7'h40),
                  $signed(reg678)}))))
            begin
              reg874 = reg709;
              reg875 <= ((reg743[(1'h1):(1'h1)] || reg720[(1'h1):(1'h0)]) != $unsigned(((~|(reg695 ?
                      reg755 : (8'ha5))) ?
                  (8'hb5) : $signed($unsigned(reg689)))));
              reg876 <= (reg761[(2'h2):(1'h1)] ?
                  (reg758[(4'hd):(2'h3)] ?
                      reg758 : (~^($signed(reg805) ^~ $signed(reg762)))) : (((wire700[(4'h8):(2'h2)] ?
                          {reg829} : $signed((8'hbf))) ?
                      ({(7'h41)} ?
                          reg820 : (~reg722)) : reg820) < wire649[(4'h8):(3'h5)]));
            end
          else
            begin
              reg875 <= $signed(((|({reg873} ?
                      (wire647 ? reg669 : reg812) : (reg791 && reg871))) ?
                  {(+(reg752 ?
                          reg876 : reg709))} : (&(reg779 && $unsigned(reg686)))));
              reg877 = (^$signed(reg657));
            end
          for (forvar878 = (1'h0); (forvar878 < (1'h0)); forvar878 = (forvar878 + (1'h1)))
            begin
              reg879 <= $unsigned(reg715[(2'h2):(1'h0)]);
              reg880 = (^$signed($unsigned((reg726[(2'h3):(2'h3)] ?
                  reg676 : wire845[(1'h1):(1'h0)]))));
            end
        end
      else
        begin
          reg874 = (!$unsigned((reg675[(3'h6):(2'h3)] ?
              ((~|reg779) ?
                  reg817[(3'h5):(3'h5)] : $signed((8'hbc))) : reg667[(2'h3):(2'h3)])));
          reg877 = reg817[(1'h1):(1'h0)];
        end
      for (forvar881 = (1'h0); (forvar881 < (2'h3)); forvar881 = (forvar881 + (1'h1)))
        begin
          if (reg869)
            begin
              reg882 = reg658;
              reg883 = {$unsigned(reg695[(2'h3):(2'h3)])};
            end
          else
            begin
              reg882 = $unsigned($signed($signed(reg723[(4'ha):(2'h3)])));
              reg883 = $signed((($unsigned((^~reg882)) ?
                      wire700 : (&(reg753 + reg754))) ?
                  $signed(((reg869 ? reg786 : wire648) ?
                      $signed(wire648) : reg686[(3'h5):(2'h2)])) : $unsigned((!$unsigned(reg807)))));
              reg884 = {$unsigned(reg810),
                  ((~&(|(reg800 ? (8'ha6) : reg675))) ?
                      (reg718[(5'h16):(4'ha)] ?
                          reg847[(3'h6):(3'h6)] : reg720[(2'h2):(1'h1)]) : $unsigned(reg712))};
              reg885 = wire648[(4'hf):(3'h7)];
              reg886 = reg785;
            end
          reg887 <= reg653;
          if ((reg718 && (^reg719)))
            begin
              reg888 = (&reg883);
              reg889 <= $unsigned(reg856);
              reg890 = $signed((8'hb0));
              reg891 <= $signed($unsigned({wire652,
                  (reg817[(4'he):(4'hd)] ~^ {reg761, reg815})}));
            end
          else
            begin
              reg889 <= $signed($signed(reg760[(3'h4):(1'h1)]));
              reg890 = ({(((~reg663) ?
                              {(8'h9d), reg792} : (reg719 ? reg695 : reg824)) ?
                          {$signed((8'ha5))} : ((~^reg737) ?
                              $signed((8'hb0)) : $unsigned(reg866)))} ?
                  ((reg829 ? {reg791, reg678} : (^(reg767 ? reg817 : reg755))) ?
                      wire647[(2'h2):(2'h2)] : reg829[(3'h4):(1'h1)]) : $unsigned((({reg876,
                          wire845} ?
                      $unsigned(reg685) : $signed(reg839)) > reg651)));
              reg892 = {((+$unsigned(wire698[(2'h3):(2'h2)])) ?
                      (~&reg806[(1'h0):(1'h0)]) : ({(reg794 == reg651)} ?
                          $signed((reg874 ?
                              (8'ha6) : (8'hbf))) : ((reg741 <= reg784) ?
                              (reg888 ? reg875 : reg847) : $signed(reg723)))),
                  ($signed(reg869) | ($signed((reg889 ? (8'ha1) : (8'hb0))) ?
                      {(+reg814)} : {reg807}))};
            end
          for (forvar893 = (1'h0); (forvar893 < (1'h0)); forvar893 = (forvar893 + (1'h1)))
            begin
              reg894 <= $signed(reg836[(1'h1):(1'h1)]);
              reg895 <= reg720[(2'h2):(1'h0)];
              reg896 = $unsigned((reg741[(1'h1):(1'h0)] ?
                  $signed($signed(reg737[(2'h2):(1'h1)])) : (reg895 ?
                      $signed((reg788 ~^ reg875)) : reg873[(5'h12):(4'h8)])));
              reg897 = reg691;
              reg898 <= reg784[(1'h1):(1'h0)];
            end
          for (forvar899 = (1'h0); (forvar899 < (2'h2)); forvar899 = (forvar899 + (1'h1)))
            begin
              reg900 <= (^($signed($unsigned((~|(8'hbe)))) == reg675[(3'h7):(2'h2)]));
              reg901 <= reg817;
              reg902 <= $signed(((|(|((7'h44) ?
                  reg812 : reg824))) >= (^reg804)));
              reg903 = (^$signed(({(reg879 & reg822)} ?
                  $signed((&reg833)) : $unsigned((^~reg762)))));
            end
        end
    end
  always
    @(posedge clk) begin
      reg904 = $signed(wire647[(3'h6):(3'h5)]);
      for (forvar905 = (1'h0); (forvar905 < (1'h1)); forvar905 = (forvar905 + (1'h1)))
        begin
          reg906 = $signed(((((wire845 == reg856) ?
                  $signed(reg725) : $unsigned(reg768)) ?
              $unsigned({reg685}) : $unsigned((~reg836))) <<< reg821));
          reg907 <= ((~&((8'hb3) >>> $unsigned($signed(reg788)))) <<< $unsigned(((~&(reg836 >= reg666)) * reg768[(5'h12):(3'h5)])));
          reg908 = $unsigned($unsigned($signed(reg786[(4'ha):(2'h2)])));
        end
      if ($unsigned(reg718[(2'h3):(1'h1)]))
        begin
          reg909 <= reg758[(4'hf):(3'h4)];
          for (forvar910 = (1'h0); (forvar910 < (2'h3)); forvar910 = (forvar910 + (1'h1)))
            begin
              reg911 = forvar905;
              reg912 <= reg821;
            end
          if ($unsigned($unsigned($signed((!(~|(8'haa)))))))
            begin
              reg913 <= ((~&(-$unsigned((reg693 ?
                  (7'h48) : reg806)))) >> reg686);
              reg914 = (((|reg807[(4'hc):(2'h3)]) ?
                      reg841 : (|{$signed(reg706)})) ?
                  reg785 : $unsigned(reg784));
              reg915 = reg894[(2'h3):(2'h3)];
            end
          else
            begin
              reg913 <= ((reg737[(1'h1):(1'h1)] ?
                  $signed($unsigned((reg712 ?
                      reg847 : reg709))) : reg833) * ($signed({(reg777 + (8'hb7)),
                      $signed(reg657)}) ?
                  reg779[(1'h0):(1'h0)] : reg814));
              reg916 <= ((!(|$unsigned((reg807 - reg765)))) ~^ $unsigned($signed(reg758[(5'h13):(4'hc)])));
            end
          reg917 = (+reg706);
        end
      else
        begin
          reg910 = $signed((wire652 ?
              $signed($signed((reg829 ?
                  reg722 : reg665))) : (($signed((8'h9d)) ?
                  (reg653 ?
                      reg760 : reg792) : $unsigned((8'hb2))) & (reg815[(4'h8):(2'h3)] ?
                  reg913[(2'h3):(1'h0)] : reg806))));
          for (forvar911 = (1'h0); (forvar911 < (2'h3)); forvar911 = (forvar911 + (1'h1)))
            begin
              reg912 <= $signed((~|reg762[(1'h1):(1'h1)]));
              reg914 = $signed((reg681 ~^ (|(reg760 ?
                  $signed(reg712) : (reg681 > reg871)))));
              reg916 <= ($signed(($unsigned($unsigned(reg853)) ?
                      $unsigned({reg715}) : $unsigned(((8'ha2) ?
                          reg807 : reg911)))) ?
                  (+$signed($unsigned(((7'h40) ? (8'hb9) : reg828)))) : reg715);
              reg917 = ({$signed(((reg666 ? reg856 : wire870) + (reg719 ?
                          reg758 : (8'h9d))))} ?
                  {reg725,
                      $unsigned($signed((reg895 == reg911)))} : ($unsigned(($signed((8'hb8)) ?
                      (reg895 <= reg693) : reg762[(2'h2):(1'h1)])) <= $signed(reg815)));
            end
          for (forvar918 = (1'h0); (forvar918 < (1'h1)); forvar918 = (forvar918 + (1'h1)))
            begin
              reg919 <= {((~$signed((reg719 ? reg725 : (8'ha3)))) ?
                      forvar911 : {({reg755} > $unsigned(reg754))})};
              reg920 = wire698;
              reg921 = reg719[(3'h4):(3'h4)];
            end
          if ((^((~&wire649) ? reg785[(4'hd):(4'h9)] : reg887)))
            begin
              reg922 <= wire647;
              reg923 <= wire647;
            end
          else
            begin
              reg922 <= $unsigned((wire646 ? reg824 : reg824[(4'hd):(2'h2)]));
              reg924 = (~|reg678[(2'h3):(1'h0)]);
              reg925 <= $signed(({(~&reg915[(1'h0):(1'h0)])} == (reg769 ?
                  $signed((reg894 ? reg817 : reg653)) : reg807)));
              reg926 = ((-reg779) == $unsigned(reg869[(3'h6):(3'h6)]));
            end
          reg927 <= (&((reg786 ?
                  $signed((reg820 ?
                      (8'haa) : wire647)) : ((reg904 != reg723) ^ reg853[(4'hd):(4'h9)])) ?
              reg723[(2'h2):(1'h1)] : ((((8'hb5) <<< reg719) >= reg806[(4'h8):(3'h4)]) ?
                  $unsigned($signed(reg738)) : $signed((7'h42)))));
        end
      reg928 <= ((&$unsigned((reg830[(5'h12):(4'hf)] < (reg737 <<< reg833)))) ?
          ($signed((7'h47)) - (~|(reg685[(5'h17):(4'ha)] >= (~&reg814)))) : $signed(reg820));
      reg929 <= {$unsigned(((~&(~|reg925)) != ($signed(wire645) == reg917[(1'h0):(1'h0)])))};
    end
  assign wire930 = ({$signed(($signed(reg895) ?
                           reg752[(2'h2):(1'h1)] : (reg790 == reg871)))} & (wire648 <<< $signed(reg741[(1'h0):(1'h0)])));
  always
    @(posedge clk) begin
      reg931 = reg767;
      reg932 <= (!$signed(((reg709 && ((8'ha4) ? reg716 : reg689)) ?
          reg812 : wire930[(5'h18):(4'hd)])));
      reg933 <= {$signed(reg898[(2'h3):(1'h1)]),
          (&({$unsigned(reg691)} || ((reg907 ? reg853 : reg925) >= reg689)))};
      for (forvar934 = (1'h0); (forvar934 < (2'h3)); forvar934 = (forvar934 + (1'h1)))
        begin
          reg935 <= $unsigned(((~$signed((~^reg820))) ?
              ($unsigned(((8'ha9) <<< wire845)) > {reg891[(4'hd):(3'h6)],
                  $signed(reg922)}) : {{$unsigned(reg670)}, (8'hbd)}));
          reg936 <= $unsigned((|(reg788[(2'h3):(2'h2)] <= ((wire930 >>> reg873) >>> $signed(reg718)))));
        end
    end
  always
    @(posedge clk) begin
      reg937 <= (!reg876[(2'h3):(1'h1)]);
      if ((&(reg769 ?
          ((+(wire700 != reg833)) >>> reg822[(3'h5):(3'h5)]) : (((|reg857) ?
                  reg829[(2'h2):(1'h1)] : (7'h46)) ?
              (~&{(8'haf)}) : ((reg810 >= reg728) ?
                  $unsigned(reg824) : (reg923 ? reg929 : reg779))))))
        begin
          if (reg719[(3'h6):(1'h1)])
            begin
              reg938 = $signed((($signed((reg810 < reg695)) ?
                      ($unsigned(reg761) ?
                          wire646 : reg866) : ((reg788 < reg687) <<< (&reg754))) ?
                  {$unsigned(reg857[(2'h2):(2'h2)])} : (-(|reg902[(4'he):(4'h9)]))));
              reg939 = $signed(reg653);
              reg940 <= ((&$signed({{reg728, (7'h4a)}})) ?
                  reg791 : (~^(reg869[(2'h2):(2'h2)] + $signed(reg839))));
              reg941 = $signed(((reg875 + ((7'h49) | {(8'ha5), reg912})) ?
                  $unsigned($signed((reg725 ? reg807 : (8'haa)))) : (8'hb7)));
            end
          else
            begin
              reg938 = wire649[(4'h9):(3'h5)];
              reg939 = reg790[(3'h5):(1'h0)];
              reg941 = ((~$unsigned((reg779 ? {reg876} : {reg676}))) ?
                  $signed(((~reg736) | reg695)) : $signed(reg847[(3'h7):(3'h7)]));
            end
          for (forvar942 = (1'h0); (forvar942 < (1'h1)); forvar942 = (forvar942 + (1'h1)))
            begin
              reg943 <= (8'ha2);
            end
          for (forvar944 = (1'h0); (forvar944 < (2'h2)); forvar944 = (forvar944 + (1'h1)))
            begin
              reg945 <= (+(~|$unsigned(((reg909 ? reg728 : reg832) >= (reg800 ?
                  wire652 : (8'ha4))))));
              reg946 = $unsigned($signed(reg714[(4'h8):(1'h0)]));
            end
        end
      else
        begin
          for (forvar938 = (1'h0); (forvar938 < (3'h4)); forvar938 = (forvar938 + (1'h1)))
            begin
              reg940 <= (($unsigned(($signed(reg933) ?
                  (|reg832) : reg788[(4'h9):(3'h5)])) | reg706) ~^ $unsigned((^~((+reg928) ?
                  (wire648 >> reg847) : reg869[(2'h3):(1'h0)]))));
              reg942 <= (~|((-((forvar942 >> reg833) ?
                  reg820[(4'ha):(2'h3)] : (reg938 ?
                      reg821 : reg737))) != {((~|reg830) && reg817)}));
              reg944 = (&reg693[(3'h6):(3'h6)]);
            end
          reg946 = $signed($signed(reg784[(3'h5):(2'h3)]));
          if ($signed(reg695[(1'h1):(1'h1)]))
            begin
              reg947 = ($unsigned((^$unsigned($signed(reg806)))) || reg682[(1'h0):(1'h0)]);
              reg948 <= $unsigned($unsigned(reg658[(3'h5):(3'h4)]));
              reg949 = reg706[(3'h7):(1'h1)];
              reg950 = ((({reg935[(3'h7):(3'h7)]} << wire845[(2'h3):(1'h0)]) & (-{(reg752 | reg871),
                      (reg907 != reg936)})) ?
                  (^$unsigned(((7'h40) ?
                      (+reg822) : $unsigned(reg919)))) : ((^~(((8'hb8) ?
                      reg682 : (7'h47)) + (8'ha6))) | (&reg754)));
              reg951 = reg857[(1'h0):(1'h0)];
            end
          else
            begin
              reg948 <= (reg789 ?
                  ($unsigned(((reg779 >= reg922) > ((8'h9e) ?
                      reg854 : reg670))) <<< ($unsigned((reg891 ?
                      reg857 : reg935)) * $signed($signed(wire870)))) : reg757);
              reg952 <= (reg792 ? (!reg830) : wire646);
              reg953 = reg932;
            end
          reg954 <= $unsigned((8'ha5));
          if ($signed((reg791 == (~|reg786))))
            begin
              reg955 <= (-({(-$signed(reg814)), $unsigned((reg820 || reg768))} ?
                  (+(7'h43)) : ((&((7'h49) ?
                      wire646 : wire844)) != (~^reg706))));
              reg956 <= (reg669[(1'h1):(1'h0)] >= (($unsigned((reg813 >> reg928)) ?
                      reg946 : (reg947[(2'h2):(1'h0)] ?
                          reg945 : reg928[(1'h0):(1'h0)])) ?
                  ($signed(reg789[(2'h2):(1'h0)]) >= {(reg869 ?
                          reg812 : reg803),
                      (reg932 ?
                          reg676 : reg762)}) : $unsigned({$unsigned(reg909),
                      reg820[(4'he):(3'h7)]})));
            end
          else
            begin
              reg955 <= {(~&reg656[(3'h4):(2'h2)]),
                  $unsigned(((7'h44) || (~^(reg654 ? reg935 : reg891))))};
              reg957 = {(($unsigned($signed(reg709)) ?
                          (reg913[(2'h3):(1'h1)] ^~ (reg752 && (7'h42))) : ((^reg715) > forvar942)) ?
                      reg901 : reg738),
                  {(8'hba), $unsigned(reg769[(5'h12):(1'h0)])}};
            end
        end
    end
  assign wire958 = reg712;
endmodule